# 
#              Synchronous High Speed Single Port SRAM Compiler 
# 
#                    UMC 0.18um GenericII Logic Process
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : SUMA180_432X44X1BM1
#       Words            : 432
#       Bits             : 44
#       Byte-Write       : 1
#       Aspect Ratio     : 1
#       Output Loading   : 0.05  (pf)
#       Data Slew        : 0.02  (ns)
#       CK Slew          : 0.02  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2024/11/03 21:47:36
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO SUMA180_432X44X1BM1
CLASS BLOCK ;
FOREIGN SUMA180_432X44X1BM1 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 726.020 BY 269.360 ;
SYMMETRY x y r90 ;
SITE core_5040 ;
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal4 ;
  RECT 724.900 255.140 726.020 258.380 ;
  LAYER metal3 ;
  RECT 724.900 255.140 726.020 258.380 ;
  LAYER metal2 ;
  RECT 724.900 255.140 726.020 258.380 ;
  LAYER metal1 ;
  RECT 724.900 255.140 726.020 258.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 247.300 726.020 250.540 ;
  LAYER metal3 ;
  RECT 724.900 247.300 726.020 250.540 ;
  LAYER metal2 ;
  RECT 724.900 247.300 726.020 250.540 ;
  LAYER metal1 ;
  RECT 724.900 247.300 726.020 250.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 208.100 726.020 211.340 ;
  LAYER metal3 ;
  RECT 724.900 208.100 726.020 211.340 ;
  LAYER metal2 ;
  RECT 724.900 208.100 726.020 211.340 ;
  LAYER metal1 ;
  RECT 724.900 208.100 726.020 211.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 200.260 726.020 203.500 ;
  LAYER metal3 ;
  RECT 724.900 200.260 726.020 203.500 ;
  LAYER metal2 ;
  RECT 724.900 200.260 726.020 203.500 ;
  LAYER metal1 ;
  RECT 724.900 200.260 726.020 203.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 192.420 726.020 195.660 ;
  LAYER metal3 ;
  RECT 724.900 192.420 726.020 195.660 ;
  LAYER metal2 ;
  RECT 724.900 192.420 726.020 195.660 ;
  LAYER metal1 ;
  RECT 724.900 192.420 726.020 195.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 184.580 726.020 187.820 ;
  LAYER metal3 ;
  RECT 724.900 184.580 726.020 187.820 ;
  LAYER metal2 ;
  RECT 724.900 184.580 726.020 187.820 ;
  LAYER metal1 ;
  RECT 724.900 184.580 726.020 187.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 176.740 726.020 179.980 ;
  LAYER metal3 ;
  RECT 724.900 176.740 726.020 179.980 ;
  LAYER metal2 ;
  RECT 724.900 176.740 726.020 179.980 ;
  LAYER metal1 ;
  RECT 724.900 176.740 726.020 179.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 168.900 726.020 172.140 ;
  LAYER metal3 ;
  RECT 724.900 168.900 726.020 172.140 ;
  LAYER metal2 ;
  RECT 724.900 168.900 726.020 172.140 ;
  LAYER metal1 ;
  RECT 724.900 168.900 726.020 172.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 129.700 726.020 132.940 ;
  LAYER metal3 ;
  RECT 724.900 129.700 726.020 132.940 ;
  LAYER metal2 ;
  RECT 724.900 129.700 726.020 132.940 ;
  LAYER metal1 ;
  RECT 724.900 129.700 726.020 132.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 121.860 726.020 125.100 ;
  LAYER metal3 ;
  RECT 724.900 121.860 726.020 125.100 ;
  LAYER metal2 ;
  RECT 724.900 121.860 726.020 125.100 ;
  LAYER metal1 ;
  RECT 724.900 121.860 726.020 125.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 114.020 726.020 117.260 ;
  LAYER metal3 ;
  RECT 724.900 114.020 726.020 117.260 ;
  LAYER metal2 ;
  RECT 724.900 114.020 726.020 117.260 ;
  LAYER metal1 ;
  RECT 724.900 114.020 726.020 117.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 106.180 726.020 109.420 ;
  LAYER metal3 ;
  RECT 724.900 106.180 726.020 109.420 ;
  LAYER metal2 ;
  RECT 724.900 106.180 726.020 109.420 ;
  LAYER metal1 ;
  RECT 724.900 106.180 726.020 109.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 98.340 726.020 101.580 ;
  LAYER metal3 ;
  RECT 724.900 98.340 726.020 101.580 ;
  LAYER metal2 ;
  RECT 724.900 98.340 726.020 101.580 ;
  LAYER metal1 ;
  RECT 724.900 98.340 726.020 101.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 90.500 726.020 93.740 ;
  LAYER metal3 ;
  RECT 724.900 90.500 726.020 93.740 ;
  LAYER metal2 ;
  RECT 724.900 90.500 726.020 93.740 ;
  LAYER metal1 ;
  RECT 724.900 90.500 726.020 93.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 51.300 726.020 54.540 ;
  LAYER metal3 ;
  RECT 724.900 51.300 726.020 54.540 ;
  LAYER metal2 ;
  RECT 724.900 51.300 726.020 54.540 ;
  LAYER metal1 ;
  RECT 724.900 51.300 726.020 54.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 43.460 726.020 46.700 ;
  LAYER metal3 ;
  RECT 724.900 43.460 726.020 46.700 ;
  LAYER metal2 ;
  RECT 724.900 43.460 726.020 46.700 ;
  LAYER metal1 ;
  RECT 724.900 43.460 726.020 46.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 35.620 726.020 38.860 ;
  LAYER metal3 ;
  RECT 724.900 35.620 726.020 38.860 ;
  LAYER metal2 ;
  RECT 724.900 35.620 726.020 38.860 ;
  LAYER metal1 ;
  RECT 724.900 35.620 726.020 38.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 27.780 726.020 31.020 ;
  LAYER metal3 ;
  RECT 724.900 27.780 726.020 31.020 ;
  LAYER metal2 ;
  RECT 724.900 27.780 726.020 31.020 ;
  LAYER metal1 ;
  RECT 724.900 27.780 726.020 31.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 19.940 726.020 23.180 ;
  LAYER metal3 ;
  RECT 724.900 19.940 726.020 23.180 ;
  LAYER metal2 ;
  RECT 724.900 19.940 726.020 23.180 ;
  LAYER metal1 ;
  RECT 724.900 19.940 726.020 23.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 12.100 726.020 15.340 ;
  LAYER metal3 ;
  RECT 724.900 12.100 726.020 15.340 ;
  LAYER metal2 ;
  RECT 724.900 12.100 726.020 15.340 ;
  LAYER metal1 ;
  RECT 724.900 12.100 726.020 15.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER metal3 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER metal2 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER metal1 ;
  RECT 0.000 255.140 1.120 258.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER metal3 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER metal2 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER metal1 ;
  RECT 0.000 247.300 1.120 250.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER metal3 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER metal2 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER metal1 ;
  RECT 0.000 208.100 1.120 211.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER metal3 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER metal2 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER metal1 ;
  RECT 0.000 200.260 1.120 203.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER metal3 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER metal2 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER metal1 ;
  RECT 0.000 192.420 1.120 195.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER metal3 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER metal2 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER metal1 ;
  RECT 0.000 184.580 1.120 187.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER metal3 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER metal2 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER metal1 ;
  RECT 0.000 176.740 1.120 179.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER metal3 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER metal2 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER metal1 ;
  RECT 0.000 168.900 1.120 172.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal3 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal2 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal1 ;
  RECT 0.000 129.700 1.120 132.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal3 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal2 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal1 ;
  RECT 0.000 121.860 1.120 125.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal3 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal2 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal1 ;
  RECT 0.000 114.020 1.120 117.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal3 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal2 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal1 ;
  RECT 0.000 106.180 1.120 109.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal3 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal2 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal1 ;
  RECT 0.000 98.340 1.120 101.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal3 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal2 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal1 ;
  RECT 0.000 90.500 1.120 93.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal3 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal2 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal1 ;
  RECT 0.000 51.300 1.120 54.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal3 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal2 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal1 ;
  RECT 0.000 43.460 1.120 46.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal3 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal2 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal1 ;
  RECT 0.000 35.620 1.120 38.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal3 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal2 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal1 ;
  RECT 0.000 27.780 1.120 31.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal3 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal2 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal1 ;
  RECT 0.000 19.940 1.120 23.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal3 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal2 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal1 ;
  RECT 0.000 12.100 1.120 15.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 706.580 268.240 710.120 269.360 ;
  LAYER metal3 ;
  RECT 706.580 268.240 710.120 269.360 ;
  LAYER metal2 ;
  RECT 706.580 268.240 710.120 269.360 ;
  LAYER metal1 ;
  RECT 706.580 268.240 710.120 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 663.180 268.240 666.720 269.360 ;
  LAYER metal3 ;
  RECT 663.180 268.240 666.720 269.360 ;
  LAYER metal2 ;
  RECT 663.180 268.240 666.720 269.360 ;
  LAYER metal1 ;
  RECT 663.180 268.240 666.720 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 654.500 268.240 658.040 269.360 ;
  LAYER metal3 ;
  RECT 654.500 268.240 658.040 269.360 ;
  LAYER metal2 ;
  RECT 654.500 268.240 658.040 269.360 ;
  LAYER metal1 ;
  RECT 654.500 268.240 658.040 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 645.820 268.240 649.360 269.360 ;
  LAYER metal3 ;
  RECT 645.820 268.240 649.360 269.360 ;
  LAYER metal2 ;
  RECT 645.820 268.240 649.360 269.360 ;
  LAYER metal1 ;
  RECT 645.820 268.240 649.360 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 637.140 268.240 640.680 269.360 ;
  LAYER metal3 ;
  RECT 637.140 268.240 640.680 269.360 ;
  LAYER metal2 ;
  RECT 637.140 268.240 640.680 269.360 ;
  LAYER metal1 ;
  RECT 637.140 268.240 640.680 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 628.460 268.240 632.000 269.360 ;
  LAYER metal3 ;
  RECT 628.460 268.240 632.000 269.360 ;
  LAYER metal2 ;
  RECT 628.460 268.240 632.000 269.360 ;
  LAYER metal1 ;
  RECT 628.460 268.240 632.000 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 619.780 268.240 623.320 269.360 ;
  LAYER metal3 ;
  RECT 619.780 268.240 623.320 269.360 ;
  LAYER metal2 ;
  RECT 619.780 268.240 623.320 269.360 ;
  LAYER metal1 ;
  RECT 619.780 268.240 623.320 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 576.380 268.240 579.920 269.360 ;
  LAYER metal3 ;
  RECT 576.380 268.240 579.920 269.360 ;
  LAYER metal2 ;
  RECT 576.380 268.240 579.920 269.360 ;
  LAYER metal1 ;
  RECT 576.380 268.240 579.920 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 567.700 268.240 571.240 269.360 ;
  LAYER metal3 ;
  RECT 567.700 268.240 571.240 269.360 ;
  LAYER metal2 ;
  RECT 567.700 268.240 571.240 269.360 ;
  LAYER metal1 ;
  RECT 567.700 268.240 571.240 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 559.020 268.240 562.560 269.360 ;
  LAYER metal3 ;
  RECT 559.020 268.240 562.560 269.360 ;
  LAYER metal2 ;
  RECT 559.020 268.240 562.560 269.360 ;
  LAYER metal1 ;
  RECT 559.020 268.240 562.560 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 550.340 268.240 553.880 269.360 ;
  LAYER metal3 ;
  RECT 550.340 268.240 553.880 269.360 ;
  LAYER metal2 ;
  RECT 550.340 268.240 553.880 269.360 ;
  LAYER metal1 ;
  RECT 550.340 268.240 553.880 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 541.660 268.240 545.200 269.360 ;
  LAYER metal3 ;
  RECT 541.660 268.240 545.200 269.360 ;
  LAYER metal2 ;
  RECT 541.660 268.240 545.200 269.360 ;
  LAYER metal1 ;
  RECT 541.660 268.240 545.200 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 532.980 268.240 536.520 269.360 ;
  LAYER metal3 ;
  RECT 532.980 268.240 536.520 269.360 ;
  LAYER metal2 ;
  RECT 532.980 268.240 536.520 269.360 ;
  LAYER metal1 ;
  RECT 532.980 268.240 536.520 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 489.580 268.240 493.120 269.360 ;
  LAYER metal3 ;
  RECT 489.580 268.240 493.120 269.360 ;
  LAYER metal2 ;
  RECT 489.580 268.240 493.120 269.360 ;
  LAYER metal1 ;
  RECT 489.580 268.240 493.120 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 480.900 268.240 484.440 269.360 ;
  LAYER metal3 ;
  RECT 480.900 268.240 484.440 269.360 ;
  LAYER metal2 ;
  RECT 480.900 268.240 484.440 269.360 ;
  LAYER metal1 ;
  RECT 480.900 268.240 484.440 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 472.220 268.240 475.760 269.360 ;
  LAYER metal3 ;
  RECT 472.220 268.240 475.760 269.360 ;
  LAYER metal2 ;
  RECT 472.220 268.240 475.760 269.360 ;
  LAYER metal1 ;
  RECT 472.220 268.240 475.760 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 463.540 268.240 467.080 269.360 ;
  LAYER metal3 ;
  RECT 463.540 268.240 467.080 269.360 ;
  LAYER metal2 ;
  RECT 463.540 268.240 467.080 269.360 ;
  LAYER metal1 ;
  RECT 463.540 268.240 467.080 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 454.860 268.240 458.400 269.360 ;
  LAYER metal3 ;
  RECT 454.860 268.240 458.400 269.360 ;
  LAYER metal2 ;
  RECT 454.860 268.240 458.400 269.360 ;
  LAYER metal1 ;
  RECT 454.860 268.240 458.400 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 446.180 268.240 449.720 269.360 ;
  LAYER metal3 ;
  RECT 446.180 268.240 449.720 269.360 ;
  LAYER metal2 ;
  RECT 446.180 268.240 449.720 269.360 ;
  LAYER metal1 ;
  RECT 446.180 268.240 449.720 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 402.780 268.240 406.320 269.360 ;
  LAYER metal3 ;
  RECT 402.780 268.240 406.320 269.360 ;
  LAYER metal2 ;
  RECT 402.780 268.240 406.320 269.360 ;
  LAYER metal1 ;
  RECT 402.780 268.240 406.320 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 394.100 268.240 397.640 269.360 ;
  LAYER metal3 ;
  RECT 394.100 268.240 397.640 269.360 ;
  LAYER metal2 ;
  RECT 394.100 268.240 397.640 269.360 ;
  LAYER metal1 ;
  RECT 394.100 268.240 397.640 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 385.420 268.240 388.960 269.360 ;
  LAYER metal3 ;
  RECT 385.420 268.240 388.960 269.360 ;
  LAYER metal2 ;
  RECT 385.420 268.240 388.960 269.360 ;
  LAYER metal1 ;
  RECT 385.420 268.240 388.960 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 376.740 268.240 380.280 269.360 ;
  LAYER metal3 ;
  RECT 376.740 268.240 380.280 269.360 ;
  LAYER metal2 ;
  RECT 376.740 268.240 380.280 269.360 ;
  LAYER metal1 ;
  RECT 376.740 268.240 380.280 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 368.060 268.240 371.600 269.360 ;
  LAYER metal3 ;
  RECT 368.060 268.240 371.600 269.360 ;
  LAYER metal2 ;
  RECT 368.060 268.240 371.600 269.360 ;
  LAYER metal1 ;
  RECT 368.060 268.240 371.600 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 359.380 268.240 362.920 269.360 ;
  LAYER metal3 ;
  RECT 359.380 268.240 362.920 269.360 ;
  LAYER metal2 ;
  RECT 359.380 268.240 362.920 269.360 ;
  LAYER metal1 ;
  RECT 359.380 268.240 362.920 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.980 268.240 319.520 269.360 ;
  LAYER metal3 ;
  RECT 315.980 268.240 319.520 269.360 ;
  LAYER metal2 ;
  RECT 315.980 268.240 319.520 269.360 ;
  LAYER metal1 ;
  RECT 315.980 268.240 319.520 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 307.300 268.240 310.840 269.360 ;
  LAYER metal3 ;
  RECT 307.300 268.240 310.840 269.360 ;
  LAYER metal2 ;
  RECT 307.300 268.240 310.840 269.360 ;
  LAYER metal1 ;
  RECT 307.300 268.240 310.840 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 298.620 268.240 302.160 269.360 ;
  LAYER metal3 ;
  RECT 298.620 268.240 302.160 269.360 ;
  LAYER metal2 ;
  RECT 298.620 268.240 302.160 269.360 ;
  LAYER metal1 ;
  RECT 298.620 268.240 302.160 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 289.940 268.240 293.480 269.360 ;
  LAYER metal3 ;
  RECT 289.940 268.240 293.480 269.360 ;
  LAYER metal2 ;
  RECT 289.940 268.240 293.480 269.360 ;
  LAYER metal1 ;
  RECT 289.940 268.240 293.480 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 281.260 268.240 284.800 269.360 ;
  LAYER metal3 ;
  RECT 281.260 268.240 284.800 269.360 ;
  LAYER metal2 ;
  RECT 281.260 268.240 284.800 269.360 ;
  LAYER metal1 ;
  RECT 281.260 268.240 284.800 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 272.580 268.240 276.120 269.360 ;
  LAYER metal3 ;
  RECT 272.580 268.240 276.120 269.360 ;
  LAYER metal2 ;
  RECT 272.580 268.240 276.120 269.360 ;
  LAYER metal1 ;
  RECT 272.580 268.240 276.120 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 229.180 268.240 232.720 269.360 ;
  LAYER metal3 ;
  RECT 229.180 268.240 232.720 269.360 ;
  LAYER metal2 ;
  RECT 229.180 268.240 232.720 269.360 ;
  LAYER metal1 ;
  RECT 229.180 268.240 232.720 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 220.500 268.240 224.040 269.360 ;
  LAYER metal3 ;
  RECT 220.500 268.240 224.040 269.360 ;
  LAYER metal2 ;
  RECT 220.500 268.240 224.040 269.360 ;
  LAYER metal1 ;
  RECT 220.500 268.240 224.040 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 211.820 268.240 215.360 269.360 ;
  LAYER metal3 ;
  RECT 211.820 268.240 215.360 269.360 ;
  LAYER metal2 ;
  RECT 211.820 268.240 215.360 269.360 ;
  LAYER metal1 ;
  RECT 211.820 268.240 215.360 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 203.140 268.240 206.680 269.360 ;
  LAYER metal3 ;
  RECT 203.140 268.240 206.680 269.360 ;
  LAYER metal2 ;
  RECT 203.140 268.240 206.680 269.360 ;
  LAYER metal1 ;
  RECT 203.140 268.240 206.680 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 194.460 268.240 198.000 269.360 ;
  LAYER metal3 ;
  RECT 194.460 268.240 198.000 269.360 ;
  LAYER metal2 ;
  RECT 194.460 268.240 198.000 269.360 ;
  LAYER metal1 ;
  RECT 194.460 268.240 198.000 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 185.780 268.240 189.320 269.360 ;
  LAYER metal3 ;
  RECT 185.780 268.240 189.320 269.360 ;
  LAYER metal2 ;
  RECT 185.780 268.240 189.320 269.360 ;
  LAYER metal1 ;
  RECT 185.780 268.240 189.320 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 142.380 268.240 145.920 269.360 ;
  LAYER metal3 ;
  RECT 142.380 268.240 145.920 269.360 ;
  LAYER metal2 ;
  RECT 142.380 268.240 145.920 269.360 ;
  LAYER metal1 ;
  RECT 142.380 268.240 145.920 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 133.700 268.240 137.240 269.360 ;
  LAYER metal3 ;
  RECT 133.700 268.240 137.240 269.360 ;
  LAYER metal2 ;
  RECT 133.700 268.240 137.240 269.360 ;
  LAYER metal1 ;
  RECT 133.700 268.240 137.240 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 125.020 268.240 128.560 269.360 ;
  LAYER metal3 ;
  RECT 125.020 268.240 128.560 269.360 ;
  LAYER metal2 ;
  RECT 125.020 268.240 128.560 269.360 ;
  LAYER metal1 ;
  RECT 125.020 268.240 128.560 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 116.340 268.240 119.880 269.360 ;
  LAYER metal3 ;
  RECT 116.340 268.240 119.880 269.360 ;
  LAYER metal2 ;
  RECT 116.340 268.240 119.880 269.360 ;
  LAYER metal1 ;
  RECT 116.340 268.240 119.880 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 107.660 268.240 111.200 269.360 ;
  LAYER metal3 ;
  RECT 107.660 268.240 111.200 269.360 ;
  LAYER metal2 ;
  RECT 107.660 268.240 111.200 269.360 ;
  LAYER metal1 ;
  RECT 107.660 268.240 111.200 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 98.980 268.240 102.520 269.360 ;
  LAYER metal3 ;
  RECT 98.980 268.240 102.520 269.360 ;
  LAYER metal2 ;
  RECT 98.980 268.240 102.520 269.360 ;
  LAYER metal1 ;
  RECT 98.980 268.240 102.520 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 55.580 268.240 59.120 269.360 ;
  LAYER metal3 ;
  RECT 55.580 268.240 59.120 269.360 ;
  LAYER metal2 ;
  RECT 55.580 268.240 59.120 269.360 ;
  LAYER metal1 ;
  RECT 55.580 268.240 59.120 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 46.900 268.240 50.440 269.360 ;
  LAYER metal3 ;
  RECT 46.900 268.240 50.440 269.360 ;
  LAYER metal2 ;
  RECT 46.900 268.240 50.440 269.360 ;
  LAYER metal1 ;
  RECT 46.900 268.240 50.440 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 38.220 268.240 41.760 269.360 ;
  LAYER metal3 ;
  RECT 38.220 268.240 41.760 269.360 ;
  LAYER metal2 ;
  RECT 38.220 268.240 41.760 269.360 ;
  LAYER metal1 ;
  RECT 38.220 268.240 41.760 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 29.540 268.240 33.080 269.360 ;
  LAYER metal3 ;
  RECT 29.540 268.240 33.080 269.360 ;
  LAYER metal2 ;
  RECT 29.540 268.240 33.080 269.360 ;
  LAYER metal1 ;
  RECT 29.540 268.240 33.080 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 20.860 268.240 24.400 269.360 ;
  LAYER metal3 ;
  RECT 20.860 268.240 24.400 269.360 ;
  LAYER metal2 ;
  RECT 20.860 268.240 24.400 269.360 ;
  LAYER metal1 ;
  RECT 20.860 268.240 24.400 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 12.180 268.240 15.720 269.360 ;
  LAYER metal3 ;
  RECT 12.180 268.240 15.720 269.360 ;
  LAYER metal2 ;
  RECT 12.180 268.240 15.720 269.360 ;
  LAYER metal1 ;
  RECT 12.180 268.240 15.720 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 714.640 0.000 718.180 1.120 ;
  LAYER metal3 ;
  RECT 714.640 0.000 718.180 1.120 ;
  LAYER metal2 ;
  RECT 714.640 0.000 718.180 1.120 ;
  LAYER metal1 ;
  RECT 714.640 0.000 718.180 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 697.900 0.000 701.440 1.120 ;
  LAYER metal3 ;
  RECT 697.900 0.000 701.440 1.120 ;
  LAYER metal2 ;
  RECT 697.900 0.000 701.440 1.120 ;
  LAYER metal1 ;
  RECT 697.900 0.000 701.440 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 676.200 0.000 679.740 1.120 ;
  LAYER metal3 ;
  RECT 676.200 0.000 679.740 1.120 ;
  LAYER metal2 ;
  RECT 676.200 0.000 679.740 1.120 ;
  LAYER metal1 ;
  RECT 676.200 0.000 679.740 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 563.360 0.000 566.900 1.120 ;
  LAYER metal3 ;
  RECT 563.360 0.000 566.900 1.120 ;
  LAYER metal2 ;
  RECT 563.360 0.000 566.900 1.120 ;
  LAYER metal1 ;
  RECT 563.360 0.000 566.900 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 541.660 0.000 545.200 1.120 ;
  LAYER metal3 ;
  RECT 541.660 0.000 545.200 1.120 ;
  LAYER metal2 ;
  RECT 541.660 0.000 545.200 1.120 ;
  LAYER metal1 ;
  RECT 541.660 0.000 545.200 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 519.960 0.000 523.500 1.120 ;
  LAYER metal3 ;
  RECT 519.960 0.000 523.500 1.120 ;
  LAYER metal2 ;
  RECT 519.960 0.000 523.500 1.120 ;
  LAYER metal1 ;
  RECT 519.960 0.000 523.500 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 493.300 0.000 496.840 1.120 ;
  LAYER metal3 ;
  RECT 493.300 0.000 496.840 1.120 ;
  LAYER metal2 ;
  RECT 493.300 0.000 496.840 1.120 ;
  LAYER metal1 ;
  RECT 493.300 0.000 496.840 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 476.560 0.000 480.100 1.120 ;
  LAYER metal3 ;
  RECT 476.560 0.000 480.100 1.120 ;
  LAYER metal2 ;
  RECT 476.560 0.000 480.100 1.120 ;
  LAYER metal1 ;
  RECT 476.560 0.000 480.100 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 449.900 0.000 453.440 1.120 ;
  LAYER metal3 ;
  RECT 449.900 0.000 453.440 1.120 ;
  LAYER metal2 ;
  RECT 449.900 0.000 453.440 1.120 ;
  LAYER metal1 ;
  RECT 449.900 0.000 453.440 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 343.260 0.000 346.800 1.120 ;
  LAYER metal3 ;
  RECT 343.260 0.000 346.800 1.120 ;
  LAYER metal2 ;
  RECT 343.260 0.000 346.800 1.120 ;
  LAYER metal1 ;
  RECT 343.260 0.000 346.800 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 325.900 0.000 329.440 1.120 ;
  LAYER metal3 ;
  RECT 325.900 0.000 329.440 1.120 ;
  LAYER metal2 ;
  RECT 325.900 0.000 329.440 1.120 ;
  LAYER metal1 ;
  RECT 325.900 0.000 329.440 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 312.880 0.000 316.420 1.120 ;
  LAYER metal3 ;
  RECT 312.880 0.000 316.420 1.120 ;
  LAYER metal2 ;
  RECT 312.880 0.000 316.420 1.120 ;
  LAYER metal1 ;
  RECT 312.880 0.000 316.420 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 296.760 0.000 300.300 1.120 ;
  LAYER metal3 ;
  RECT 296.760 0.000 300.300 1.120 ;
  LAYER metal2 ;
  RECT 296.760 0.000 300.300 1.120 ;
  LAYER metal1 ;
  RECT 296.760 0.000 300.300 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 270.100 0.000 273.640 1.120 ;
  LAYER metal3 ;
  RECT 270.100 0.000 273.640 1.120 ;
  LAYER metal2 ;
  RECT 270.100 0.000 273.640 1.120 ;
  LAYER metal1 ;
  RECT 270.100 0.000 273.640 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER metal3 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER metal2 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER metal1 ;
  RECT 253.360 0.000 256.900 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER metal3 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER metal2 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER metal1 ;
  RECT 139.900 0.000 143.440 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER metal3 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER metal2 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER metal1 ;
  RECT 113.860 0.000 117.400 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER metal3 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER metal2 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER metal1 ;
  RECT 92.160 0.000 95.700 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal3 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal2 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal1 ;
  RECT 70.460 0.000 74.000 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER metal3 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER metal2 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER metal1 ;
  RECT 43.800 0.000 47.340 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal3 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal2 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal1 ;
  RECT 27.060 0.000 30.600 1.120 ;
 END
END GND
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal4 ;
  RECT 724.900 251.220 726.020 254.460 ;
  LAYER metal3 ;
  RECT 724.900 251.220 726.020 254.460 ;
  LAYER metal2 ;
  RECT 724.900 251.220 726.020 254.460 ;
  LAYER metal1 ;
  RECT 724.900 251.220 726.020 254.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 243.380 726.020 246.620 ;
  LAYER metal3 ;
  RECT 724.900 243.380 726.020 246.620 ;
  LAYER metal2 ;
  RECT 724.900 243.380 726.020 246.620 ;
  LAYER metal1 ;
  RECT 724.900 243.380 726.020 246.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 204.180 726.020 207.420 ;
  LAYER metal3 ;
  RECT 724.900 204.180 726.020 207.420 ;
  LAYER metal2 ;
  RECT 724.900 204.180 726.020 207.420 ;
  LAYER metal1 ;
  RECT 724.900 204.180 726.020 207.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 196.340 726.020 199.580 ;
  LAYER metal3 ;
  RECT 724.900 196.340 726.020 199.580 ;
  LAYER metal2 ;
  RECT 724.900 196.340 726.020 199.580 ;
  LAYER metal1 ;
  RECT 724.900 196.340 726.020 199.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 188.500 726.020 191.740 ;
  LAYER metal3 ;
  RECT 724.900 188.500 726.020 191.740 ;
  LAYER metal2 ;
  RECT 724.900 188.500 726.020 191.740 ;
  LAYER metal1 ;
  RECT 724.900 188.500 726.020 191.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 180.660 726.020 183.900 ;
  LAYER metal3 ;
  RECT 724.900 180.660 726.020 183.900 ;
  LAYER metal2 ;
  RECT 724.900 180.660 726.020 183.900 ;
  LAYER metal1 ;
  RECT 724.900 180.660 726.020 183.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 172.820 726.020 176.060 ;
  LAYER metal3 ;
  RECT 724.900 172.820 726.020 176.060 ;
  LAYER metal2 ;
  RECT 724.900 172.820 726.020 176.060 ;
  LAYER metal1 ;
  RECT 724.900 172.820 726.020 176.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 164.980 726.020 168.220 ;
  LAYER metal3 ;
  RECT 724.900 164.980 726.020 168.220 ;
  LAYER metal2 ;
  RECT 724.900 164.980 726.020 168.220 ;
  LAYER metal1 ;
  RECT 724.900 164.980 726.020 168.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 125.780 726.020 129.020 ;
  LAYER metal3 ;
  RECT 724.900 125.780 726.020 129.020 ;
  LAYER metal2 ;
  RECT 724.900 125.780 726.020 129.020 ;
  LAYER metal1 ;
  RECT 724.900 125.780 726.020 129.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 117.940 726.020 121.180 ;
  LAYER metal3 ;
  RECT 724.900 117.940 726.020 121.180 ;
  LAYER metal2 ;
  RECT 724.900 117.940 726.020 121.180 ;
  LAYER metal1 ;
  RECT 724.900 117.940 726.020 121.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 110.100 726.020 113.340 ;
  LAYER metal3 ;
  RECT 724.900 110.100 726.020 113.340 ;
  LAYER metal2 ;
  RECT 724.900 110.100 726.020 113.340 ;
  LAYER metal1 ;
  RECT 724.900 110.100 726.020 113.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 102.260 726.020 105.500 ;
  LAYER metal3 ;
  RECT 724.900 102.260 726.020 105.500 ;
  LAYER metal2 ;
  RECT 724.900 102.260 726.020 105.500 ;
  LAYER metal1 ;
  RECT 724.900 102.260 726.020 105.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 94.420 726.020 97.660 ;
  LAYER metal3 ;
  RECT 724.900 94.420 726.020 97.660 ;
  LAYER metal2 ;
  RECT 724.900 94.420 726.020 97.660 ;
  LAYER metal1 ;
  RECT 724.900 94.420 726.020 97.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 86.580 726.020 89.820 ;
  LAYER metal3 ;
  RECT 724.900 86.580 726.020 89.820 ;
  LAYER metal2 ;
  RECT 724.900 86.580 726.020 89.820 ;
  LAYER metal1 ;
  RECT 724.900 86.580 726.020 89.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 47.380 726.020 50.620 ;
  LAYER metal3 ;
  RECT 724.900 47.380 726.020 50.620 ;
  LAYER metal2 ;
  RECT 724.900 47.380 726.020 50.620 ;
  LAYER metal1 ;
  RECT 724.900 47.380 726.020 50.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 39.540 726.020 42.780 ;
  LAYER metal3 ;
  RECT 724.900 39.540 726.020 42.780 ;
  LAYER metal2 ;
  RECT 724.900 39.540 726.020 42.780 ;
  LAYER metal1 ;
  RECT 724.900 39.540 726.020 42.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 31.700 726.020 34.940 ;
  LAYER metal3 ;
  RECT 724.900 31.700 726.020 34.940 ;
  LAYER metal2 ;
  RECT 724.900 31.700 726.020 34.940 ;
  LAYER metal1 ;
  RECT 724.900 31.700 726.020 34.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 23.860 726.020 27.100 ;
  LAYER metal3 ;
  RECT 724.900 23.860 726.020 27.100 ;
  LAYER metal2 ;
  RECT 724.900 23.860 726.020 27.100 ;
  LAYER metal1 ;
  RECT 724.900 23.860 726.020 27.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 16.020 726.020 19.260 ;
  LAYER metal3 ;
  RECT 724.900 16.020 726.020 19.260 ;
  LAYER metal2 ;
  RECT 724.900 16.020 726.020 19.260 ;
  LAYER metal1 ;
  RECT 724.900 16.020 726.020 19.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 724.900 8.180 726.020 11.420 ;
  LAYER metal3 ;
  RECT 724.900 8.180 726.020 11.420 ;
  LAYER metal2 ;
  RECT 724.900 8.180 726.020 11.420 ;
  LAYER metal1 ;
  RECT 724.900 8.180 726.020 11.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER metal3 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER metal2 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER metal1 ;
  RECT 0.000 251.220 1.120 254.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER metal3 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER metal2 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER metal1 ;
  RECT 0.000 243.380 1.120 246.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER metal3 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER metal2 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER metal1 ;
  RECT 0.000 204.180 1.120 207.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER metal3 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER metal2 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER metal1 ;
  RECT 0.000 196.340 1.120 199.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER metal3 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER metal2 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER metal1 ;
  RECT 0.000 188.500 1.120 191.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER metal3 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER metal2 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER metal1 ;
  RECT 0.000 180.660 1.120 183.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER metal3 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER metal2 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER metal1 ;
  RECT 0.000 172.820 1.120 176.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER metal3 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER metal2 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER metal1 ;
  RECT 0.000 164.980 1.120 168.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal3 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal2 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal1 ;
  RECT 0.000 125.780 1.120 129.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal3 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal2 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal1 ;
  RECT 0.000 117.940 1.120 121.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal3 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal2 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal1 ;
  RECT 0.000 110.100 1.120 113.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal3 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal2 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal1 ;
  RECT 0.000 102.260 1.120 105.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal3 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal2 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal1 ;
  RECT 0.000 94.420 1.120 97.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal3 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal2 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal1 ;
  RECT 0.000 86.580 1.120 89.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal3 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal2 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal1 ;
  RECT 0.000 47.380 1.120 50.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal3 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal2 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal1 ;
  RECT 0.000 39.540 1.120 42.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal3 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal2 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal1 ;
  RECT 0.000 31.700 1.120 34.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal3 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal2 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal1 ;
  RECT 0.000 23.860 1.120 27.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal3 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal2 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal1 ;
  RECT 0.000 16.020 1.120 19.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal3 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal2 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal1 ;
  RECT 0.000 8.180 1.120 11.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 710.920 268.240 714.460 269.360 ;
  LAYER metal3 ;
  RECT 710.920 268.240 714.460 269.360 ;
  LAYER metal2 ;
  RECT 710.920 268.240 714.460 269.360 ;
  LAYER metal1 ;
  RECT 710.920 268.240 714.460 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 702.240 268.240 705.780 269.360 ;
  LAYER metal3 ;
  RECT 702.240 268.240 705.780 269.360 ;
  LAYER metal2 ;
  RECT 702.240 268.240 705.780 269.360 ;
  LAYER metal1 ;
  RECT 702.240 268.240 705.780 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 658.840 268.240 662.380 269.360 ;
  LAYER metal3 ;
  RECT 658.840 268.240 662.380 269.360 ;
  LAYER metal2 ;
  RECT 658.840 268.240 662.380 269.360 ;
  LAYER metal1 ;
  RECT 658.840 268.240 662.380 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 650.160 268.240 653.700 269.360 ;
  LAYER metal3 ;
  RECT 650.160 268.240 653.700 269.360 ;
  LAYER metal2 ;
  RECT 650.160 268.240 653.700 269.360 ;
  LAYER metal1 ;
  RECT 650.160 268.240 653.700 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 641.480 268.240 645.020 269.360 ;
  LAYER metal3 ;
  RECT 641.480 268.240 645.020 269.360 ;
  LAYER metal2 ;
  RECT 641.480 268.240 645.020 269.360 ;
  LAYER metal1 ;
  RECT 641.480 268.240 645.020 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 632.800 268.240 636.340 269.360 ;
  LAYER metal3 ;
  RECT 632.800 268.240 636.340 269.360 ;
  LAYER metal2 ;
  RECT 632.800 268.240 636.340 269.360 ;
  LAYER metal1 ;
  RECT 632.800 268.240 636.340 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 624.120 268.240 627.660 269.360 ;
  LAYER metal3 ;
  RECT 624.120 268.240 627.660 269.360 ;
  LAYER metal2 ;
  RECT 624.120 268.240 627.660 269.360 ;
  LAYER metal1 ;
  RECT 624.120 268.240 627.660 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 615.440 268.240 618.980 269.360 ;
  LAYER metal3 ;
  RECT 615.440 268.240 618.980 269.360 ;
  LAYER metal2 ;
  RECT 615.440 268.240 618.980 269.360 ;
  LAYER metal1 ;
  RECT 615.440 268.240 618.980 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 572.040 268.240 575.580 269.360 ;
  LAYER metal3 ;
  RECT 572.040 268.240 575.580 269.360 ;
  LAYER metal2 ;
  RECT 572.040 268.240 575.580 269.360 ;
  LAYER metal1 ;
  RECT 572.040 268.240 575.580 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 563.360 268.240 566.900 269.360 ;
  LAYER metal3 ;
  RECT 563.360 268.240 566.900 269.360 ;
  LAYER metal2 ;
  RECT 563.360 268.240 566.900 269.360 ;
  LAYER metal1 ;
  RECT 563.360 268.240 566.900 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 554.680 268.240 558.220 269.360 ;
  LAYER metal3 ;
  RECT 554.680 268.240 558.220 269.360 ;
  LAYER metal2 ;
  RECT 554.680 268.240 558.220 269.360 ;
  LAYER metal1 ;
  RECT 554.680 268.240 558.220 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 546.000 268.240 549.540 269.360 ;
  LAYER metal3 ;
  RECT 546.000 268.240 549.540 269.360 ;
  LAYER metal2 ;
  RECT 546.000 268.240 549.540 269.360 ;
  LAYER metal1 ;
  RECT 546.000 268.240 549.540 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 537.320 268.240 540.860 269.360 ;
  LAYER metal3 ;
  RECT 537.320 268.240 540.860 269.360 ;
  LAYER metal2 ;
  RECT 537.320 268.240 540.860 269.360 ;
  LAYER metal1 ;
  RECT 537.320 268.240 540.860 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 528.640 268.240 532.180 269.360 ;
  LAYER metal3 ;
  RECT 528.640 268.240 532.180 269.360 ;
  LAYER metal2 ;
  RECT 528.640 268.240 532.180 269.360 ;
  LAYER metal1 ;
  RECT 528.640 268.240 532.180 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 485.240 268.240 488.780 269.360 ;
  LAYER metal3 ;
  RECT 485.240 268.240 488.780 269.360 ;
  LAYER metal2 ;
  RECT 485.240 268.240 488.780 269.360 ;
  LAYER metal1 ;
  RECT 485.240 268.240 488.780 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 476.560 268.240 480.100 269.360 ;
  LAYER metal3 ;
  RECT 476.560 268.240 480.100 269.360 ;
  LAYER metal2 ;
  RECT 476.560 268.240 480.100 269.360 ;
  LAYER metal1 ;
  RECT 476.560 268.240 480.100 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 467.880 268.240 471.420 269.360 ;
  LAYER metal3 ;
  RECT 467.880 268.240 471.420 269.360 ;
  LAYER metal2 ;
  RECT 467.880 268.240 471.420 269.360 ;
  LAYER metal1 ;
  RECT 467.880 268.240 471.420 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 459.200 268.240 462.740 269.360 ;
  LAYER metal3 ;
  RECT 459.200 268.240 462.740 269.360 ;
  LAYER metal2 ;
  RECT 459.200 268.240 462.740 269.360 ;
  LAYER metal1 ;
  RECT 459.200 268.240 462.740 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 450.520 268.240 454.060 269.360 ;
  LAYER metal3 ;
  RECT 450.520 268.240 454.060 269.360 ;
  LAYER metal2 ;
  RECT 450.520 268.240 454.060 269.360 ;
  LAYER metal1 ;
  RECT 450.520 268.240 454.060 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 441.840 268.240 445.380 269.360 ;
  LAYER metal3 ;
  RECT 441.840 268.240 445.380 269.360 ;
  LAYER metal2 ;
  RECT 441.840 268.240 445.380 269.360 ;
  LAYER metal1 ;
  RECT 441.840 268.240 445.380 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 398.440 268.240 401.980 269.360 ;
  LAYER metal3 ;
  RECT 398.440 268.240 401.980 269.360 ;
  LAYER metal2 ;
  RECT 398.440 268.240 401.980 269.360 ;
  LAYER metal1 ;
  RECT 398.440 268.240 401.980 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 389.760 268.240 393.300 269.360 ;
  LAYER metal3 ;
  RECT 389.760 268.240 393.300 269.360 ;
  LAYER metal2 ;
  RECT 389.760 268.240 393.300 269.360 ;
  LAYER metal1 ;
  RECT 389.760 268.240 393.300 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 381.080 268.240 384.620 269.360 ;
  LAYER metal3 ;
  RECT 381.080 268.240 384.620 269.360 ;
  LAYER metal2 ;
  RECT 381.080 268.240 384.620 269.360 ;
  LAYER metal1 ;
  RECT 381.080 268.240 384.620 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 372.400 268.240 375.940 269.360 ;
  LAYER metal3 ;
  RECT 372.400 268.240 375.940 269.360 ;
  LAYER metal2 ;
  RECT 372.400 268.240 375.940 269.360 ;
  LAYER metal1 ;
  RECT 372.400 268.240 375.940 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 363.720 268.240 367.260 269.360 ;
  LAYER metal3 ;
  RECT 363.720 268.240 367.260 269.360 ;
  LAYER metal2 ;
  RECT 363.720 268.240 367.260 269.360 ;
  LAYER metal1 ;
  RECT 363.720 268.240 367.260 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 355.040 268.240 358.580 269.360 ;
  LAYER metal3 ;
  RECT 355.040 268.240 358.580 269.360 ;
  LAYER metal2 ;
  RECT 355.040 268.240 358.580 269.360 ;
  LAYER metal1 ;
  RECT 355.040 268.240 358.580 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 311.640 268.240 315.180 269.360 ;
  LAYER metal3 ;
  RECT 311.640 268.240 315.180 269.360 ;
  LAYER metal2 ;
  RECT 311.640 268.240 315.180 269.360 ;
  LAYER metal1 ;
  RECT 311.640 268.240 315.180 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 302.960 268.240 306.500 269.360 ;
  LAYER metal3 ;
  RECT 302.960 268.240 306.500 269.360 ;
  LAYER metal2 ;
  RECT 302.960 268.240 306.500 269.360 ;
  LAYER metal1 ;
  RECT 302.960 268.240 306.500 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 294.280 268.240 297.820 269.360 ;
  LAYER metal3 ;
  RECT 294.280 268.240 297.820 269.360 ;
  LAYER metal2 ;
  RECT 294.280 268.240 297.820 269.360 ;
  LAYER metal1 ;
  RECT 294.280 268.240 297.820 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 285.600 268.240 289.140 269.360 ;
  LAYER metal3 ;
  RECT 285.600 268.240 289.140 269.360 ;
  LAYER metal2 ;
  RECT 285.600 268.240 289.140 269.360 ;
  LAYER metal1 ;
  RECT 285.600 268.240 289.140 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 276.920 268.240 280.460 269.360 ;
  LAYER metal3 ;
  RECT 276.920 268.240 280.460 269.360 ;
  LAYER metal2 ;
  RECT 276.920 268.240 280.460 269.360 ;
  LAYER metal1 ;
  RECT 276.920 268.240 280.460 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 268.240 268.240 271.780 269.360 ;
  LAYER metal3 ;
  RECT 268.240 268.240 271.780 269.360 ;
  LAYER metal2 ;
  RECT 268.240 268.240 271.780 269.360 ;
  LAYER metal1 ;
  RECT 268.240 268.240 271.780 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 224.840 268.240 228.380 269.360 ;
  LAYER metal3 ;
  RECT 224.840 268.240 228.380 269.360 ;
  LAYER metal2 ;
  RECT 224.840 268.240 228.380 269.360 ;
  LAYER metal1 ;
  RECT 224.840 268.240 228.380 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 216.160 268.240 219.700 269.360 ;
  LAYER metal3 ;
  RECT 216.160 268.240 219.700 269.360 ;
  LAYER metal2 ;
  RECT 216.160 268.240 219.700 269.360 ;
  LAYER metal1 ;
  RECT 216.160 268.240 219.700 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 207.480 268.240 211.020 269.360 ;
  LAYER metal3 ;
  RECT 207.480 268.240 211.020 269.360 ;
  LAYER metal2 ;
  RECT 207.480 268.240 211.020 269.360 ;
  LAYER metal1 ;
  RECT 207.480 268.240 211.020 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 198.800 268.240 202.340 269.360 ;
  LAYER metal3 ;
  RECT 198.800 268.240 202.340 269.360 ;
  LAYER metal2 ;
  RECT 198.800 268.240 202.340 269.360 ;
  LAYER metal1 ;
  RECT 198.800 268.240 202.340 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 190.120 268.240 193.660 269.360 ;
  LAYER metal3 ;
  RECT 190.120 268.240 193.660 269.360 ;
  LAYER metal2 ;
  RECT 190.120 268.240 193.660 269.360 ;
  LAYER metal1 ;
  RECT 190.120 268.240 193.660 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 181.440 268.240 184.980 269.360 ;
  LAYER metal3 ;
  RECT 181.440 268.240 184.980 269.360 ;
  LAYER metal2 ;
  RECT 181.440 268.240 184.980 269.360 ;
  LAYER metal1 ;
  RECT 181.440 268.240 184.980 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 138.040 268.240 141.580 269.360 ;
  LAYER metal3 ;
  RECT 138.040 268.240 141.580 269.360 ;
  LAYER metal2 ;
  RECT 138.040 268.240 141.580 269.360 ;
  LAYER metal1 ;
  RECT 138.040 268.240 141.580 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 129.360 268.240 132.900 269.360 ;
  LAYER metal3 ;
  RECT 129.360 268.240 132.900 269.360 ;
  LAYER metal2 ;
  RECT 129.360 268.240 132.900 269.360 ;
  LAYER metal1 ;
  RECT 129.360 268.240 132.900 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 120.680 268.240 124.220 269.360 ;
  LAYER metal3 ;
  RECT 120.680 268.240 124.220 269.360 ;
  LAYER metal2 ;
  RECT 120.680 268.240 124.220 269.360 ;
  LAYER metal1 ;
  RECT 120.680 268.240 124.220 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 112.000 268.240 115.540 269.360 ;
  LAYER metal3 ;
  RECT 112.000 268.240 115.540 269.360 ;
  LAYER metal2 ;
  RECT 112.000 268.240 115.540 269.360 ;
  LAYER metal1 ;
  RECT 112.000 268.240 115.540 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 103.320 268.240 106.860 269.360 ;
  LAYER metal3 ;
  RECT 103.320 268.240 106.860 269.360 ;
  LAYER metal2 ;
  RECT 103.320 268.240 106.860 269.360 ;
  LAYER metal1 ;
  RECT 103.320 268.240 106.860 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 94.640 268.240 98.180 269.360 ;
  LAYER metal3 ;
  RECT 94.640 268.240 98.180 269.360 ;
  LAYER metal2 ;
  RECT 94.640 268.240 98.180 269.360 ;
  LAYER metal1 ;
  RECT 94.640 268.240 98.180 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 51.240 268.240 54.780 269.360 ;
  LAYER metal3 ;
  RECT 51.240 268.240 54.780 269.360 ;
  LAYER metal2 ;
  RECT 51.240 268.240 54.780 269.360 ;
  LAYER metal1 ;
  RECT 51.240 268.240 54.780 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 42.560 268.240 46.100 269.360 ;
  LAYER metal3 ;
  RECT 42.560 268.240 46.100 269.360 ;
  LAYER metal2 ;
  RECT 42.560 268.240 46.100 269.360 ;
  LAYER metal1 ;
  RECT 42.560 268.240 46.100 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 33.880 268.240 37.420 269.360 ;
  LAYER metal3 ;
  RECT 33.880 268.240 37.420 269.360 ;
  LAYER metal2 ;
  RECT 33.880 268.240 37.420 269.360 ;
  LAYER metal1 ;
  RECT 33.880 268.240 37.420 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 25.200 268.240 28.740 269.360 ;
  LAYER metal3 ;
  RECT 25.200 268.240 28.740 269.360 ;
  LAYER metal2 ;
  RECT 25.200 268.240 28.740 269.360 ;
  LAYER metal1 ;
  RECT 25.200 268.240 28.740 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 16.520 268.240 20.060 269.360 ;
  LAYER metal3 ;
  RECT 16.520 268.240 20.060 269.360 ;
  LAYER metal2 ;
  RECT 16.520 268.240 20.060 269.360 ;
  LAYER metal1 ;
  RECT 16.520 268.240 20.060 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 7.840 268.240 11.380 269.360 ;
  LAYER metal3 ;
  RECT 7.840 268.240 11.380 269.360 ;
  LAYER metal2 ;
  RECT 7.840 268.240 11.380 269.360 ;
  LAYER metal1 ;
  RECT 7.840 268.240 11.380 269.360 ;
 END
 PORT
  LAYER metal4 ;
  RECT 705.960 0.000 709.500 1.120 ;
  LAYER metal3 ;
  RECT 705.960 0.000 709.500 1.120 ;
  LAYER metal2 ;
  RECT 705.960 0.000 709.500 1.120 ;
  LAYER metal1 ;
  RECT 705.960 0.000 709.500 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 689.220 0.000 692.760 1.120 ;
  LAYER metal3 ;
  RECT 689.220 0.000 692.760 1.120 ;
  LAYER metal2 ;
  RECT 689.220 0.000 692.760 1.120 ;
  LAYER metal1 ;
  RECT 689.220 0.000 692.760 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 663.180 0.000 666.720 1.120 ;
  LAYER metal3 ;
  RECT 663.180 0.000 666.720 1.120 ;
  LAYER metal2 ;
  RECT 663.180 0.000 666.720 1.120 ;
  LAYER metal1 ;
  RECT 663.180 0.000 666.720 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 549.720 0.000 553.260 1.120 ;
  LAYER metal3 ;
  RECT 549.720 0.000 553.260 1.120 ;
  LAYER metal2 ;
  RECT 549.720 0.000 553.260 1.120 ;
  LAYER metal1 ;
  RECT 549.720 0.000 553.260 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 532.980 0.000 536.520 1.120 ;
  LAYER metal3 ;
  RECT 532.980 0.000 536.520 1.120 ;
  LAYER metal2 ;
  RECT 532.980 0.000 536.520 1.120 ;
  LAYER metal1 ;
  RECT 532.980 0.000 536.520 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 506.940 0.000 510.480 1.120 ;
  LAYER metal3 ;
  RECT 506.940 0.000 510.480 1.120 ;
  LAYER metal2 ;
  RECT 506.940 0.000 510.480 1.120 ;
  LAYER metal1 ;
  RECT 506.940 0.000 510.480 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 485.240 0.000 488.780 1.120 ;
  LAYER metal3 ;
  RECT 485.240 0.000 488.780 1.120 ;
  LAYER metal2 ;
  RECT 485.240 0.000 488.780 1.120 ;
  LAYER metal1 ;
  RECT 485.240 0.000 488.780 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 463.540 0.000 467.080 1.120 ;
  LAYER metal3 ;
  RECT 463.540 0.000 467.080 1.120 ;
  LAYER metal2 ;
  RECT 463.540 0.000 467.080 1.120 ;
  LAYER metal1 ;
  RECT 463.540 0.000 467.080 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 436.880 0.000 440.420 1.120 ;
  LAYER metal3 ;
  RECT 436.880 0.000 440.420 1.120 ;
  LAYER metal2 ;
  RECT 436.880 0.000 440.420 1.120 ;
  LAYER metal1 ;
  RECT 436.880 0.000 440.420 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 332.720 0.000 336.260 1.120 ;
  LAYER metal3 ;
  RECT 332.720 0.000 336.260 1.120 ;
  LAYER metal2 ;
  RECT 332.720 0.000 336.260 1.120 ;
  LAYER metal1 ;
  RECT 332.720 0.000 336.260 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 321.560 0.000 325.100 1.120 ;
  LAYER metal3 ;
  RECT 321.560 0.000 325.100 1.120 ;
  LAYER metal2 ;
  RECT 321.560 0.000 325.100 1.120 ;
  LAYER metal1 ;
  RECT 321.560 0.000 325.100 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 304.820 0.000 308.360 1.120 ;
  LAYER metal3 ;
  RECT 304.820 0.000 308.360 1.120 ;
  LAYER metal2 ;
  RECT 304.820 0.000 308.360 1.120 ;
  LAYER metal1 ;
  RECT 304.820 0.000 308.360 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER metal3 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER metal2 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER metal1 ;
  RECT 283.120 0.000 286.660 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER metal3 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER metal2 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER metal1 ;
  RECT 261.420 0.000 264.960 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER metal3 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER metal2 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER metal1 ;
  RECT 239.720 0.000 243.260 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER metal3 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER metal2 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER metal1 ;
  RECT 126.880 0.000 130.420 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER metal3 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER metal2 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER metal1 ;
  RECT 100.220 0.000 103.760 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER metal3 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER metal2 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER metal1 ;
  RECT 83.480 0.000 87.020 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER metal3 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER metal2 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER metal1 ;
  RECT 56.820 0.000 60.360 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal3 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal2 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal1 ;
  RECT 35.740 0.000 39.280 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal3 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal2 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal1 ;
  RECT 14.040 0.000 17.580 1.120 ;
 END
END VCC
PIN DO43
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 712.440 0.000 713.560 1.120 ;
  LAYER metal3 ;
  RECT 712.440 0.000 713.560 1.120 ;
  LAYER metal2 ;
  RECT 712.440 0.000 713.560 1.120 ;
  LAYER metal1 ;
  RECT 712.440 0.000 713.560 1.120 ;
 END
END DO43
PIN DI43
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 703.760 0.000 704.880 1.120 ;
  LAYER metal3 ;
  RECT 703.760 0.000 704.880 1.120 ;
  LAYER metal2 ;
  RECT 703.760 0.000 704.880 1.120 ;
  LAYER metal1 ;
  RECT 703.760 0.000 704.880 1.120 ;
 END
END DI43
PIN DO42
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 695.700 0.000 696.820 1.120 ;
  LAYER metal3 ;
  RECT 695.700 0.000 696.820 1.120 ;
  LAYER metal2 ;
  RECT 695.700 0.000 696.820 1.120 ;
  LAYER metal1 ;
  RECT 695.700 0.000 696.820 1.120 ;
 END
END DO42
PIN DI42
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 687.020 0.000 688.140 1.120 ;
  LAYER metal3 ;
  RECT 687.020 0.000 688.140 1.120 ;
  LAYER metal2 ;
  RECT 687.020 0.000 688.140 1.120 ;
  LAYER metal1 ;
  RECT 687.020 0.000 688.140 1.120 ;
 END
END DI42
PIN DO41
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 682.680 0.000 683.800 1.120 ;
  LAYER metal3 ;
  RECT 682.680 0.000 683.800 1.120 ;
  LAYER metal2 ;
  RECT 682.680 0.000 683.800 1.120 ;
  LAYER metal1 ;
  RECT 682.680 0.000 683.800 1.120 ;
 END
END DO41
PIN DI41
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 674.000 0.000 675.120 1.120 ;
  LAYER metal3 ;
  RECT 674.000 0.000 675.120 1.120 ;
  LAYER metal2 ;
  RECT 674.000 0.000 675.120 1.120 ;
  LAYER metal1 ;
  RECT 674.000 0.000 675.120 1.120 ;
 END
END DI41
PIN DO40
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 669.040 0.000 670.160 1.120 ;
  LAYER metal3 ;
  RECT 669.040 0.000 670.160 1.120 ;
  LAYER metal2 ;
  RECT 669.040 0.000 670.160 1.120 ;
  LAYER metal1 ;
  RECT 669.040 0.000 670.160 1.120 ;
 END
END DO40
PIN DI40
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 660.980 0.000 662.100 1.120 ;
  LAYER metal3 ;
  RECT 660.980 0.000 662.100 1.120 ;
  LAYER metal2 ;
  RECT 660.980 0.000 662.100 1.120 ;
  LAYER metal1 ;
  RECT 660.980 0.000 662.100 1.120 ;
 END
END DI40
PIN DO39
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 652.300 0.000 653.420 1.120 ;
  LAYER metal3 ;
  RECT 652.300 0.000 653.420 1.120 ;
  LAYER metal2 ;
  RECT 652.300 0.000 653.420 1.120 ;
  LAYER metal1 ;
  RECT 652.300 0.000 653.420 1.120 ;
 END
END DO39
PIN DI39
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 644.240 0.000 645.360 1.120 ;
  LAYER metal3 ;
  RECT 644.240 0.000 645.360 1.120 ;
  LAYER metal2 ;
  RECT 644.240 0.000 645.360 1.120 ;
  LAYER metal1 ;
  RECT 644.240 0.000 645.360 1.120 ;
 END
END DI39
PIN DO38
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 639.280 0.000 640.400 1.120 ;
  LAYER metal3 ;
  RECT 639.280 0.000 640.400 1.120 ;
  LAYER metal2 ;
  RECT 639.280 0.000 640.400 1.120 ;
  LAYER metal1 ;
  RECT 639.280 0.000 640.400 1.120 ;
 END
END DO38
PIN DI38
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 630.600 0.000 631.720 1.120 ;
  LAYER metal3 ;
  RECT 630.600 0.000 631.720 1.120 ;
  LAYER metal2 ;
  RECT 630.600 0.000 631.720 1.120 ;
  LAYER metal1 ;
  RECT 630.600 0.000 631.720 1.120 ;
 END
END DI38
PIN DO37
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 625.640 0.000 626.760 1.120 ;
  LAYER metal3 ;
  RECT 625.640 0.000 626.760 1.120 ;
  LAYER metal2 ;
  RECT 625.640 0.000 626.760 1.120 ;
  LAYER metal1 ;
  RECT 625.640 0.000 626.760 1.120 ;
 END
END DO37
PIN DI37
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 617.580 0.000 618.700 1.120 ;
  LAYER metal3 ;
  RECT 617.580 0.000 618.700 1.120 ;
  LAYER metal2 ;
  RECT 617.580 0.000 618.700 1.120 ;
  LAYER metal1 ;
  RECT 617.580 0.000 618.700 1.120 ;
 END
END DI37
PIN DO36
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 612.620 0.000 613.740 1.120 ;
  LAYER metal3 ;
  RECT 612.620 0.000 613.740 1.120 ;
  LAYER metal2 ;
  RECT 612.620 0.000 613.740 1.120 ;
  LAYER metal1 ;
  RECT 612.620 0.000 613.740 1.120 ;
 END
END DO36
PIN DI36
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 603.940 0.000 605.060 1.120 ;
  LAYER metal3 ;
  RECT 603.940 0.000 605.060 1.120 ;
  LAYER metal2 ;
  RECT 603.940 0.000 605.060 1.120 ;
  LAYER metal1 ;
  RECT 603.940 0.000 605.060 1.120 ;
 END
END DI36
PIN DO35
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 595.880 0.000 597.000 1.120 ;
  LAYER metal3 ;
  RECT 595.880 0.000 597.000 1.120 ;
  LAYER metal2 ;
  RECT 595.880 0.000 597.000 1.120 ;
  LAYER metal1 ;
  RECT 595.880 0.000 597.000 1.120 ;
 END
END DO35
PIN DI35
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 587.820 0.000 588.940 1.120 ;
  LAYER metal3 ;
  RECT 587.820 0.000 588.940 1.120 ;
  LAYER metal2 ;
  RECT 587.820 0.000 588.940 1.120 ;
  LAYER metal1 ;
  RECT 587.820 0.000 588.940 1.120 ;
 END
END DI35
PIN DO34
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 582.860 0.000 583.980 1.120 ;
  LAYER metal3 ;
  RECT 582.860 0.000 583.980 1.120 ;
  LAYER metal2 ;
  RECT 582.860 0.000 583.980 1.120 ;
  LAYER metal1 ;
  RECT 582.860 0.000 583.980 1.120 ;
 END
END DO34
PIN DI34
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 574.180 0.000 575.300 1.120 ;
  LAYER metal3 ;
  RECT 574.180 0.000 575.300 1.120 ;
  LAYER metal2 ;
  RECT 574.180 0.000 575.300 1.120 ;
  LAYER metal1 ;
  RECT 574.180 0.000 575.300 1.120 ;
 END
END DI34
PIN DO33
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 569.220 0.000 570.340 1.120 ;
  LAYER metal3 ;
  RECT 569.220 0.000 570.340 1.120 ;
  LAYER metal2 ;
  RECT 569.220 0.000 570.340 1.120 ;
  LAYER metal1 ;
  RECT 569.220 0.000 570.340 1.120 ;
 END
END DO33
PIN DI33
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 561.160 0.000 562.280 1.120 ;
  LAYER metal3 ;
  RECT 561.160 0.000 562.280 1.120 ;
  LAYER metal2 ;
  RECT 561.160 0.000 562.280 1.120 ;
  LAYER metal1 ;
  RECT 561.160 0.000 562.280 1.120 ;
 END
END DI33
PIN DO32
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 556.200 0.000 557.320 1.120 ;
  LAYER metal3 ;
  RECT 556.200 0.000 557.320 1.120 ;
  LAYER metal2 ;
  RECT 556.200 0.000 557.320 1.120 ;
  LAYER metal1 ;
  RECT 556.200 0.000 557.320 1.120 ;
 END
END DO32
PIN DI32
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 547.520 0.000 548.640 1.120 ;
  LAYER metal3 ;
  RECT 547.520 0.000 548.640 1.120 ;
  LAYER metal2 ;
  RECT 547.520 0.000 548.640 1.120 ;
  LAYER metal1 ;
  RECT 547.520 0.000 548.640 1.120 ;
 END
END DI32
PIN DO31
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 539.460 0.000 540.580 1.120 ;
  LAYER metal3 ;
  RECT 539.460 0.000 540.580 1.120 ;
  LAYER metal2 ;
  RECT 539.460 0.000 540.580 1.120 ;
  LAYER metal1 ;
  RECT 539.460 0.000 540.580 1.120 ;
 END
END DO31
PIN DI31
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 530.780 0.000 531.900 1.120 ;
  LAYER metal3 ;
  RECT 530.780 0.000 531.900 1.120 ;
  LAYER metal2 ;
  RECT 530.780 0.000 531.900 1.120 ;
  LAYER metal1 ;
  RECT 530.780 0.000 531.900 1.120 ;
 END
END DI31
PIN DO30
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 525.820 0.000 526.940 1.120 ;
  LAYER metal3 ;
  RECT 525.820 0.000 526.940 1.120 ;
  LAYER metal2 ;
  RECT 525.820 0.000 526.940 1.120 ;
  LAYER metal1 ;
  RECT 525.820 0.000 526.940 1.120 ;
 END
END DO30
PIN DI30
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 517.760 0.000 518.880 1.120 ;
  LAYER metal3 ;
  RECT 517.760 0.000 518.880 1.120 ;
  LAYER metal2 ;
  RECT 517.760 0.000 518.880 1.120 ;
  LAYER metal1 ;
  RECT 517.760 0.000 518.880 1.120 ;
 END
END DI30
PIN DO29
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 512.800 0.000 513.920 1.120 ;
  LAYER metal3 ;
  RECT 512.800 0.000 513.920 1.120 ;
  LAYER metal2 ;
  RECT 512.800 0.000 513.920 1.120 ;
  LAYER metal1 ;
  RECT 512.800 0.000 513.920 1.120 ;
 END
END DO29
PIN DI29
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 504.740 0.000 505.860 1.120 ;
  LAYER metal3 ;
  RECT 504.740 0.000 505.860 1.120 ;
  LAYER metal2 ;
  RECT 504.740 0.000 505.860 1.120 ;
  LAYER metal1 ;
  RECT 504.740 0.000 505.860 1.120 ;
 END
END DI29
PIN DO28
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 499.780 0.000 500.900 1.120 ;
  LAYER metal3 ;
  RECT 499.780 0.000 500.900 1.120 ;
  LAYER metal2 ;
  RECT 499.780 0.000 500.900 1.120 ;
  LAYER metal1 ;
  RECT 499.780 0.000 500.900 1.120 ;
 END
END DO28
PIN DI28
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 491.100 0.000 492.220 1.120 ;
  LAYER metal3 ;
  RECT 491.100 0.000 492.220 1.120 ;
  LAYER metal2 ;
  RECT 491.100 0.000 492.220 1.120 ;
  LAYER metal1 ;
  RECT 491.100 0.000 492.220 1.120 ;
 END
END DI28
PIN DO27
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 483.040 0.000 484.160 1.120 ;
  LAYER metal3 ;
  RECT 483.040 0.000 484.160 1.120 ;
  LAYER metal2 ;
  RECT 483.040 0.000 484.160 1.120 ;
  LAYER metal1 ;
  RECT 483.040 0.000 484.160 1.120 ;
 END
END DO27
PIN DI27
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 474.360 0.000 475.480 1.120 ;
  LAYER metal3 ;
  RECT 474.360 0.000 475.480 1.120 ;
  LAYER metal2 ;
  RECT 474.360 0.000 475.480 1.120 ;
  LAYER metal1 ;
  RECT 474.360 0.000 475.480 1.120 ;
 END
END DI27
PIN DO26
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 469.400 0.000 470.520 1.120 ;
  LAYER metal3 ;
  RECT 469.400 0.000 470.520 1.120 ;
  LAYER metal2 ;
  RECT 469.400 0.000 470.520 1.120 ;
  LAYER metal1 ;
  RECT 469.400 0.000 470.520 1.120 ;
 END
END DO26
PIN DI26
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 461.340 0.000 462.460 1.120 ;
  LAYER metal3 ;
  RECT 461.340 0.000 462.460 1.120 ;
  LAYER metal2 ;
  RECT 461.340 0.000 462.460 1.120 ;
  LAYER metal1 ;
  RECT 461.340 0.000 462.460 1.120 ;
 END
END DI26
PIN DO25
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 456.380 0.000 457.500 1.120 ;
  LAYER metal3 ;
  RECT 456.380 0.000 457.500 1.120 ;
  LAYER metal2 ;
  RECT 456.380 0.000 457.500 1.120 ;
  LAYER metal1 ;
  RECT 456.380 0.000 457.500 1.120 ;
 END
END DO25
PIN DI25
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 447.700 0.000 448.820 1.120 ;
  LAYER metal3 ;
  RECT 447.700 0.000 448.820 1.120 ;
  LAYER metal2 ;
  RECT 447.700 0.000 448.820 1.120 ;
  LAYER metal1 ;
  RECT 447.700 0.000 448.820 1.120 ;
 END
END DI25
PIN DO24
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 442.740 0.000 443.860 1.120 ;
  LAYER metal3 ;
  RECT 442.740 0.000 443.860 1.120 ;
  LAYER metal2 ;
  RECT 442.740 0.000 443.860 1.120 ;
  LAYER metal1 ;
  RECT 442.740 0.000 443.860 1.120 ;
 END
END DO24
PIN DI24
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 434.680 0.000 435.800 1.120 ;
  LAYER metal3 ;
  RECT 434.680 0.000 435.800 1.120 ;
  LAYER metal2 ;
  RECT 434.680 0.000 435.800 1.120 ;
  LAYER metal1 ;
  RECT 434.680 0.000 435.800 1.120 ;
 END
END DI24
PIN DO23
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 426.620 0.000 427.740 1.120 ;
  LAYER metal3 ;
  RECT 426.620 0.000 427.740 1.120 ;
  LAYER metal2 ;
  RECT 426.620 0.000 427.740 1.120 ;
  LAYER metal1 ;
  RECT 426.620 0.000 427.740 1.120 ;
 END
END DO23
PIN DI23
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 417.940 0.000 419.060 1.120 ;
  LAYER metal3 ;
  RECT 417.940 0.000 419.060 1.120 ;
  LAYER metal2 ;
  RECT 417.940 0.000 419.060 1.120 ;
  LAYER metal1 ;
  RECT 417.940 0.000 419.060 1.120 ;
 END
END DI23
PIN DO22
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 412.980 0.000 414.100 1.120 ;
  LAYER metal3 ;
  RECT 412.980 0.000 414.100 1.120 ;
  LAYER metal2 ;
  RECT 412.980 0.000 414.100 1.120 ;
  LAYER metal1 ;
  RECT 412.980 0.000 414.100 1.120 ;
 END
END DO22
PIN DI22
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 404.920 0.000 406.040 1.120 ;
  LAYER metal3 ;
  RECT 404.920 0.000 406.040 1.120 ;
  LAYER metal2 ;
  RECT 404.920 0.000 406.040 1.120 ;
  LAYER metal1 ;
  RECT 404.920 0.000 406.040 1.120 ;
 END
END DI22
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 399.340 0.000 400.460 1.120 ;
  LAYER metal3 ;
  RECT 399.340 0.000 400.460 1.120 ;
  LAYER metal2 ;
  RECT 399.340 0.000 400.460 1.120 ;
  LAYER metal1 ;
  RECT 399.340 0.000 400.460 1.120 ;
 END
END A1
PIN WEB
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 397.480 0.000 398.600 1.120 ;
  LAYER metal3 ;
  RECT 397.480 0.000 398.600 1.120 ;
  LAYER metal2 ;
  RECT 397.480 0.000 398.600 1.120 ;
  LAYER metal1 ;
  RECT 397.480 0.000 398.600 1.120 ;
 END
END WEB
PIN OE
  DIRECTION INPUT ;
  CAPACITANCE 0.033 ;
 PORT
  LAYER metal4 ;
  RECT 392.520 0.000 393.640 1.120 ;
  LAYER metal3 ;
  RECT 392.520 0.000 393.640 1.120 ;
  LAYER metal2 ;
  RECT 392.520 0.000 393.640 1.120 ;
  LAYER metal1 ;
  RECT 392.520 0.000 393.640 1.120 ;
 END
END OE
PIN CS
  DIRECTION INPUT ;
  CAPACITANCE 0.123 ;
 PORT
  LAYER metal4 ;
  RECT 390.660 0.000 391.780 1.120 ;
  LAYER metal3 ;
  RECT 390.660 0.000 391.780 1.120 ;
  LAYER metal2 ;
  RECT 390.660 0.000 391.780 1.120 ;
  LAYER metal1 ;
  RECT 390.660 0.000 391.780 1.120 ;
 END
END CS
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 368.960 0.000 370.080 1.120 ;
  LAYER metal3 ;
  RECT 368.960 0.000 370.080 1.120 ;
  LAYER metal2 ;
  RECT 368.960 0.000 370.080 1.120 ;
  LAYER metal1 ;
  RECT 368.960 0.000 370.080 1.120 ;
 END
END A2
PIN CK
  DIRECTION INPUT ;
  CAPACITANCE 0.063 ;
 PORT
  LAYER metal4 ;
  RECT 365.860 0.000 366.980 1.120 ;
  LAYER metal3 ;
  RECT 365.860 0.000 366.980 1.120 ;
  LAYER metal2 ;
  RECT 365.860 0.000 366.980 1.120 ;
  LAYER metal1 ;
  RECT 365.860 0.000 366.980 1.120 ;
 END
END CK
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 363.380 0.000 364.500 1.120 ;
  LAYER metal3 ;
  RECT 363.380 0.000 364.500 1.120 ;
  LAYER metal2 ;
  RECT 363.380 0.000 364.500 1.120 ;
  LAYER metal1 ;
  RECT 363.380 0.000 364.500 1.120 ;
 END
END A0
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER metal3 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER metal2 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER metal1 ;
  RECT 359.040 0.000 360.160 1.120 ;
 END
END A3
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 351.600 0.000 352.720 1.120 ;
  LAYER metal3 ;
  RECT 351.600 0.000 352.720 1.120 ;
  LAYER metal2 ;
  RECT 351.600 0.000 352.720 1.120 ;
  LAYER metal1 ;
  RECT 351.600 0.000 352.720 1.120 ;
 END
END A4
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER metal3 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER metal2 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER metal1 ;
  RECT 348.500 0.000 349.620 1.120 ;
 END
END A5
PIN A6
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 341.060 0.000 342.180 1.120 ;
  LAYER metal3 ;
  RECT 341.060 0.000 342.180 1.120 ;
  LAYER metal2 ;
  RECT 341.060 0.000 342.180 1.120 ;
  LAYER metal1 ;
  RECT 341.060 0.000 342.180 1.120 ;
 END
END A6
PIN A7
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 337.960 0.000 339.080 1.120 ;
  LAYER metal3 ;
  RECT 337.960 0.000 339.080 1.120 ;
  LAYER metal2 ;
  RECT 337.960 0.000 339.080 1.120 ;
  LAYER metal1 ;
  RECT 337.960 0.000 339.080 1.120 ;
 END
END A7
PIN A8
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 330.520 0.000 331.640 1.120 ;
  LAYER metal3 ;
  RECT 330.520 0.000 331.640 1.120 ;
  LAYER metal2 ;
  RECT 330.520 0.000 331.640 1.120 ;
  LAYER metal1 ;
  RECT 330.520 0.000 331.640 1.120 ;
 END
END A8
PIN DO21
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 319.360 0.000 320.480 1.120 ;
  LAYER metal3 ;
  RECT 319.360 0.000 320.480 1.120 ;
  LAYER metal2 ;
  RECT 319.360 0.000 320.480 1.120 ;
  LAYER metal1 ;
  RECT 319.360 0.000 320.480 1.120 ;
 END
END DO21
PIN DI21
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 310.680 0.000 311.800 1.120 ;
  LAYER metal3 ;
  RECT 310.680 0.000 311.800 1.120 ;
  LAYER metal2 ;
  RECT 310.680 0.000 311.800 1.120 ;
  LAYER metal1 ;
  RECT 310.680 0.000 311.800 1.120 ;
 END
END DI21
PIN DO20
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 302.620 0.000 303.740 1.120 ;
  LAYER metal3 ;
  RECT 302.620 0.000 303.740 1.120 ;
  LAYER metal2 ;
  RECT 302.620 0.000 303.740 1.120 ;
  LAYER metal1 ;
  RECT 302.620 0.000 303.740 1.120 ;
 END
END DO20
PIN DI20
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 294.560 0.000 295.680 1.120 ;
  LAYER metal3 ;
  RECT 294.560 0.000 295.680 1.120 ;
  LAYER metal2 ;
  RECT 294.560 0.000 295.680 1.120 ;
  LAYER metal1 ;
  RECT 294.560 0.000 295.680 1.120 ;
 END
END DI20
PIN DO19
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 289.600 0.000 290.720 1.120 ;
  LAYER metal3 ;
  RECT 289.600 0.000 290.720 1.120 ;
  LAYER metal2 ;
  RECT 289.600 0.000 290.720 1.120 ;
  LAYER metal1 ;
  RECT 289.600 0.000 290.720 1.120 ;
 END
END DO19
PIN DI19
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 280.920 0.000 282.040 1.120 ;
  LAYER metal3 ;
  RECT 280.920 0.000 282.040 1.120 ;
  LAYER metal2 ;
  RECT 280.920 0.000 282.040 1.120 ;
  LAYER metal1 ;
  RECT 280.920 0.000 282.040 1.120 ;
 END
END DI19
PIN DO18
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 275.960 0.000 277.080 1.120 ;
  LAYER metal3 ;
  RECT 275.960 0.000 277.080 1.120 ;
  LAYER metal2 ;
  RECT 275.960 0.000 277.080 1.120 ;
  LAYER metal1 ;
  RECT 275.960 0.000 277.080 1.120 ;
 END
END DO18
PIN DI18
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal3 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal2 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal1 ;
  RECT 267.900 0.000 269.020 1.120 ;
 END
END DI18
PIN DO17
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER metal3 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER metal2 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER metal1 ;
  RECT 259.220 0.000 260.340 1.120 ;
 END
END DO17
PIN DI17
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER metal3 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER metal2 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER metal1 ;
  RECT 251.160 0.000 252.280 1.120 ;
 END
END DI17
PIN DO16
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER metal3 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER metal2 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER metal1 ;
  RECT 246.200 0.000 247.320 1.120 ;
 END
END DO16
PIN DI16
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER metal3 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER metal2 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER metal1 ;
  RECT 237.520 0.000 238.640 1.120 ;
 END
END DI16
PIN DO15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER metal3 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER metal2 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER metal1 ;
  RECT 233.180 0.000 234.300 1.120 ;
 END
END DO15
PIN DI15
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER metal3 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER metal2 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER metal1 ;
  RECT 224.500 0.000 225.620 1.120 ;
 END
END DI15
PIN DO14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER metal3 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER metal2 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER metal1 ;
  RECT 219.540 0.000 220.660 1.120 ;
 END
END DO14
PIN DI14
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER metal3 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER metal2 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER metal1 ;
  RECT 211.480 0.000 212.600 1.120 ;
 END
END DI14
PIN DO13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER metal3 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER metal2 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER metal1 ;
  RECT 202.800 0.000 203.920 1.120 ;
 END
END DO13
PIN DI13
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER metal3 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER metal2 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER metal1 ;
  RECT 194.740 0.000 195.860 1.120 ;
 END
END DI13
PIN DO12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER metal3 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER metal2 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER metal1 ;
  RECT 189.780 0.000 190.900 1.120 ;
 END
END DO12
PIN DI12
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER metal3 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER metal2 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER metal1 ;
  RECT 181.100 0.000 182.220 1.120 ;
 END
END DI12
PIN DO11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER metal3 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER metal2 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER metal1 ;
  RECT 176.140 0.000 177.260 1.120 ;
 END
END DO11
PIN DI11
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER metal3 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER metal2 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER metal1 ;
  RECT 168.080 0.000 169.200 1.120 ;
 END
END DI11
PIN DO10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER metal3 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER metal2 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER metal1 ;
  RECT 163.120 0.000 164.240 1.120 ;
 END
END DO10
PIN DI10
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER metal3 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER metal2 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER metal1 ;
  RECT 154.440 0.000 155.560 1.120 ;
 END
END DI10
PIN DO9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER metal3 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER metal2 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER metal1 ;
  RECT 146.380 0.000 147.500 1.120 ;
 END
END DO9
PIN DI9
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER metal3 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER metal2 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER metal1 ;
  RECT 137.700 0.000 138.820 1.120 ;
 END
END DI9
PIN DO8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER metal3 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER metal2 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER metal1 ;
  RECT 133.360 0.000 134.480 1.120 ;
 END
END DO8
PIN DI8
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER metal3 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER metal2 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER metal1 ;
  RECT 124.680 0.000 125.800 1.120 ;
 END
END DI8
PIN DO7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER metal3 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER metal2 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER metal1 ;
  RECT 119.720 0.000 120.840 1.120 ;
 END
END DO7
PIN DI7
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER metal3 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER metal2 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER metal1 ;
  RECT 111.660 0.000 112.780 1.120 ;
 END
END DI7
PIN DO6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal3 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal2 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal1 ;
  RECT 106.700 0.000 107.820 1.120 ;
 END
END DO6
PIN DI6
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER metal3 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER metal2 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER metal1 ;
  RECT 98.020 0.000 99.140 1.120 ;
 END
END DI6
PIN DO5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER metal3 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER metal2 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER metal1 ;
  RECT 89.960 0.000 91.080 1.120 ;
 END
END DO5
PIN DI5
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER metal3 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER metal2 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER metal1 ;
  RECT 81.280 0.000 82.400 1.120 ;
 END
END DI5
PIN DO4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER metal3 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER metal2 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER metal1 ;
  RECT 76.320 0.000 77.440 1.120 ;
 END
END DO4
PIN DI4
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER metal3 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER metal2 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER metal1 ;
  RECT 68.260 0.000 69.380 1.120 ;
 END
END DI4
PIN DO3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER metal3 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER metal2 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER metal1 ;
  RECT 63.300 0.000 64.420 1.120 ;
 END
END DO3
PIN DI3
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER metal3 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER metal2 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER metal1 ;
  RECT 54.620 0.000 55.740 1.120 ;
 END
END DI3
PIN DO2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER metal3 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER metal2 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER metal1 ;
  RECT 50.280 0.000 51.400 1.120 ;
 END
END DO2
PIN DI2
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER metal3 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER metal2 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER metal1 ;
  RECT 41.600 0.000 42.720 1.120 ;
 END
END DI2
PIN DO1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal3 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal2 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal1 ;
  RECT 33.540 0.000 34.660 1.120 ;
 END
END DO1
PIN DI1
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal3 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal2 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal1 ;
  RECT 24.860 0.000 25.980 1.120 ;
 END
END DI1
PIN DO0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal3 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal2 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal1 ;
  RECT 19.900 0.000 21.020 1.120 ;
 END
END DO0
PIN DI0
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal3 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal2 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal1 ;
  RECT 11.840 0.000 12.960 1.120 ;
 END
END DI0
OBS
  LAYER metal1 SPACING 0.280 ;
  RECT 0.000 0.140 726.020 269.360 ;
  LAYER metal2 SPACING 0.320 ;
  RECT 0.000 0.140 726.020 269.360 ;
  LAYER metal3 SPACING 0.320 ;
  RECT 0.000 0.140 726.020 269.360 ;
  LAYER metal4 SPACING 0.600 ;
  RECT 0.000 0.140 726.020 269.360 ;
  LAYER via ;
  RECT 0.000 0.140 726.020 269.360 ;
  LAYER via2 ;
  RECT 0.000 0.140 726.020 269.360 ;
  LAYER via3 ;
  RECT 0.000 0.140 726.020 269.360 ;
END
END SUMA180_432X44X1BM1
END LIBRARY



