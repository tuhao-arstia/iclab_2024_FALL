# 
#              Synchronous High Speed Single Port SRAM Compiler 
# 
#                    UMC 0.18um GenericII Logic Process
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : SUMA180_288X48X1BM1
#       Words            : 288
#       Bits             : 48
#       Byte-Write       : 1
#       Aspect Ratio     : 1
#       Output Loading   : 0.05  (pf)
#       Data Slew        : 0.02  (ns)
#       CK Slew          : 0.02  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2024/11/01 22:42:24
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO SUMA180_288X48X1BM1
CLASS BLOCK ;
FOREIGN SUMA180_288X48X1BM1 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 778.720 BY 225.680 ;
SYMMETRY x y r90 ;
SITE core_5040 ;
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal4 ;
  RECT 777.600 208.100 778.720 211.340 ;
  LAYER metal3 ;
  RECT 777.600 208.100 778.720 211.340 ;
  LAYER metal2 ;
  RECT 777.600 208.100 778.720 211.340 ;
  LAYER metal1 ;
  RECT 777.600 208.100 778.720 211.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 200.260 778.720 203.500 ;
  LAYER metal3 ;
  RECT 777.600 200.260 778.720 203.500 ;
  LAYER metal2 ;
  RECT 777.600 200.260 778.720 203.500 ;
  LAYER metal1 ;
  RECT 777.600 200.260 778.720 203.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 192.420 778.720 195.660 ;
  LAYER metal3 ;
  RECT 777.600 192.420 778.720 195.660 ;
  LAYER metal2 ;
  RECT 777.600 192.420 778.720 195.660 ;
  LAYER metal1 ;
  RECT 777.600 192.420 778.720 195.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 184.580 778.720 187.820 ;
  LAYER metal3 ;
  RECT 777.600 184.580 778.720 187.820 ;
  LAYER metal2 ;
  RECT 777.600 184.580 778.720 187.820 ;
  LAYER metal1 ;
  RECT 777.600 184.580 778.720 187.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 176.740 778.720 179.980 ;
  LAYER metal3 ;
  RECT 777.600 176.740 778.720 179.980 ;
  LAYER metal2 ;
  RECT 777.600 176.740 778.720 179.980 ;
  LAYER metal1 ;
  RECT 777.600 176.740 778.720 179.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 168.900 778.720 172.140 ;
  LAYER metal3 ;
  RECT 777.600 168.900 778.720 172.140 ;
  LAYER metal2 ;
  RECT 777.600 168.900 778.720 172.140 ;
  LAYER metal1 ;
  RECT 777.600 168.900 778.720 172.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 129.700 778.720 132.940 ;
  LAYER metal3 ;
  RECT 777.600 129.700 778.720 132.940 ;
  LAYER metal2 ;
  RECT 777.600 129.700 778.720 132.940 ;
  LAYER metal1 ;
  RECT 777.600 129.700 778.720 132.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 121.860 778.720 125.100 ;
  LAYER metal3 ;
  RECT 777.600 121.860 778.720 125.100 ;
  LAYER metal2 ;
  RECT 777.600 121.860 778.720 125.100 ;
  LAYER metal1 ;
  RECT 777.600 121.860 778.720 125.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 114.020 778.720 117.260 ;
  LAYER metal3 ;
  RECT 777.600 114.020 778.720 117.260 ;
  LAYER metal2 ;
  RECT 777.600 114.020 778.720 117.260 ;
  LAYER metal1 ;
  RECT 777.600 114.020 778.720 117.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 106.180 778.720 109.420 ;
  LAYER metal3 ;
  RECT 777.600 106.180 778.720 109.420 ;
  LAYER metal2 ;
  RECT 777.600 106.180 778.720 109.420 ;
  LAYER metal1 ;
  RECT 777.600 106.180 778.720 109.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 98.340 778.720 101.580 ;
  LAYER metal3 ;
  RECT 777.600 98.340 778.720 101.580 ;
  LAYER metal2 ;
  RECT 777.600 98.340 778.720 101.580 ;
  LAYER metal1 ;
  RECT 777.600 98.340 778.720 101.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 90.500 778.720 93.740 ;
  LAYER metal3 ;
  RECT 777.600 90.500 778.720 93.740 ;
  LAYER metal2 ;
  RECT 777.600 90.500 778.720 93.740 ;
  LAYER metal1 ;
  RECT 777.600 90.500 778.720 93.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 51.300 778.720 54.540 ;
  LAYER metal3 ;
  RECT 777.600 51.300 778.720 54.540 ;
  LAYER metal2 ;
  RECT 777.600 51.300 778.720 54.540 ;
  LAYER metal1 ;
  RECT 777.600 51.300 778.720 54.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 43.460 778.720 46.700 ;
  LAYER metal3 ;
  RECT 777.600 43.460 778.720 46.700 ;
  LAYER metal2 ;
  RECT 777.600 43.460 778.720 46.700 ;
  LAYER metal1 ;
  RECT 777.600 43.460 778.720 46.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 35.620 778.720 38.860 ;
  LAYER metal3 ;
  RECT 777.600 35.620 778.720 38.860 ;
  LAYER metal2 ;
  RECT 777.600 35.620 778.720 38.860 ;
  LAYER metal1 ;
  RECT 777.600 35.620 778.720 38.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 27.780 778.720 31.020 ;
  LAYER metal3 ;
  RECT 777.600 27.780 778.720 31.020 ;
  LAYER metal2 ;
  RECT 777.600 27.780 778.720 31.020 ;
  LAYER metal1 ;
  RECT 777.600 27.780 778.720 31.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 19.940 778.720 23.180 ;
  LAYER metal3 ;
  RECT 777.600 19.940 778.720 23.180 ;
  LAYER metal2 ;
  RECT 777.600 19.940 778.720 23.180 ;
  LAYER metal1 ;
  RECT 777.600 19.940 778.720 23.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 12.100 778.720 15.340 ;
  LAYER metal3 ;
  RECT 777.600 12.100 778.720 15.340 ;
  LAYER metal2 ;
  RECT 777.600 12.100 778.720 15.340 ;
  LAYER metal1 ;
  RECT 777.600 12.100 778.720 15.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER metal3 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER metal2 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER metal1 ;
  RECT 0.000 208.100 1.120 211.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER metal3 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER metal2 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER metal1 ;
  RECT 0.000 200.260 1.120 203.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER metal3 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER metal2 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER metal1 ;
  RECT 0.000 192.420 1.120 195.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER metal3 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER metal2 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER metal1 ;
  RECT 0.000 184.580 1.120 187.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER metal3 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER metal2 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER metal1 ;
  RECT 0.000 176.740 1.120 179.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER metal3 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER metal2 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER metal1 ;
  RECT 0.000 168.900 1.120 172.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal3 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal2 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal1 ;
  RECT 0.000 129.700 1.120 132.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal3 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal2 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal1 ;
  RECT 0.000 121.860 1.120 125.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal3 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal2 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal1 ;
  RECT 0.000 114.020 1.120 117.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal3 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal2 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal1 ;
  RECT 0.000 106.180 1.120 109.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal3 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal2 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal1 ;
  RECT 0.000 98.340 1.120 101.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal3 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal2 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal1 ;
  RECT 0.000 90.500 1.120 93.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal3 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal2 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal1 ;
  RECT 0.000 51.300 1.120 54.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal3 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal2 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal1 ;
  RECT 0.000 43.460 1.120 46.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal3 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal2 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal1 ;
  RECT 0.000 35.620 1.120 38.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal3 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal2 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal1 ;
  RECT 0.000 27.780 1.120 31.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal3 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal2 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal1 ;
  RECT 0.000 19.940 1.120 23.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal3 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal2 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal1 ;
  RECT 0.000 12.100 1.120 15.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 749.980 224.560 753.520 225.680 ;
  LAYER metal3 ;
  RECT 749.980 224.560 753.520 225.680 ;
  LAYER metal2 ;
  RECT 749.980 224.560 753.520 225.680 ;
  LAYER metal1 ;
  RECT 749.980 224.560 753.520 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 741.300 224.560 744.840 225.680 ;
  LAYER metal3 ;
  RECT 741.300 224.560 744.840 225.680 ;
  LAYER metal2 ;
  RECT 741.300 224.560 744.840 225.680 ;
  LAYER metal1 ;
  RECT 741.300 224.560 744.840 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 732.620 224.560 736.160 225.680 ;
  LAYER metal3 ;
  RECT 732.620 224.560 736.160 225.680 ;
  LAYER metal2 ;
  RECT 732.620 224.560 736.160 225.680 ;
  LAYER metal1 ;
  RECT 732.620 224.560 736.160 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 723.940 224.560 727.480 225.680 ;
  LAYER metal3 ;
  RECT 723.940 224.560 727.480 225.680 ;
  LAYER metal2 ;
  RECT 723.940 224.560 727.480 225.680 ;
  LAYER metal1 ;
  RECT 723.940 224.560 727.480 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 715.260 224.560 718.800 225.680 ;
  LAYER metal3 ;
  RECT 715.260 224.560 718.800 225.680 ;
  LAYER metal2 ;
  RECT 715.260 224.560 718.800 225.680 ;
  LAYER metal1 ;
  RECT 715.260 224.560 718.800 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 706.580 224.560 710.120 225.680 ;
  LAYER metal3 ;
  RECT 706.580 224.560 710.120 225.680 ;
  LAYER metal2 ;
  RECT 706.580 224.560 710.120 225.680 ;
  LAYER metal1 ;
  RECT 706.580 224.560 710.120 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 663.180 224.560 666.720 225.680 ;
  LAYER metal3 ;
  RECT 663.180 224.560 666.720 225.680 ;
  LAYER metal2 ;
  RECT 663.180 224.560 666.720 225.680 ;
  LAYER metal1 ;
  RECT 663.180 224.560 666.720 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 654.500 224.560 658.040 225.680 ;
  LAYER metal3 ;
  RECT 654.500 224.560 658.040 225.680 ;
  LAYER metal2 ;
  RECT 654.500 224.560 658.040 225.680 ;
  LAYER metal1 ;
  RECT 654.500 224.560 658.040 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 645.820 224.560 649.360 225.680 ;
  LAYER metal3 ;
  RECT 645.820 224.560 649.360 225.680 ;
  LAYER metal2 ;
  RECT 645.820 224.560 649.360 225.680 ;
  LAYER metal1 ;
  RECT 645.820 224.560 649.360 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 637.140 224.560 640.680 225.680 ;
  LAYER metal3 ;
  RECT 637.140 224.560 640.680 225.680 ;
  LAYER metal2 ;
  RECT 637.140 224.560 640.680 225.680 ;
  LAYER metal1 ;
  RECT 637.140 224.560 640.680 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 628.460 224.560 632.000 225.680 ;
  LAYER metal3 ;
  RECT 628.460 224.560 632.000 225.680 ;
  LAYER metal2 ;
  RECT 628.460 224.560 632.000 225.680 ;
  LAYER metal1 ;
  RECT 628.460 224.560 632.000 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 619.780 224.560 623.320 225.680 ;
  LAYER metal3 ;
  RECT 619.780 224.560 623.320 225.680 ;
  LAYER metal2 ;
  RECT 619.780 224.560 623.320 225.680 ;
  LAYER metal1 ;
  RECT 619.780 224.560 623.320 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 576.380 224.560 579.920 225.680 ;
  LAYER metal3 ;
  RECT 576.380 224.560 579.920 225.680 ;
  LAYER metal2 ;
  RECT 576.380 224.560 579.920 225.680 ;
  LAYER metal1 ;
  RECT 576.380 224.560 579.920 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 567.700 224.560 571.240 225.680 ;
  LAYER metal3 ;
  RECT 567.700 224.560 571.240 225.680 ;
  LAYER metal2 ;
  RECT 567.700 224.560 571.240 225.680 ;
  LAYER metal1 ;
  RECT 567.700 224.560 571.240 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 559.020 224.560 562.560 225.680 ;
  LAYER metal3 ;
  RECT 559.020 224.560 562.560 225.680 ;
  LAYER metal2 ;
  RECT 559.020 224.560 562.560 225.680 ;
  LAYER metal1 ;
  RECT 559.020 224.560 562.560 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 550.340 224.560 553.880 225.680 ;
  LAYER metal3 ;
  RECT 550.340 224.560 553.880 225.680 ;
  LAYER metal2 ;
  RECT 550.340 224.560 553.880 225.680 ;
  LAYER metal1 ;
  RECT 550.340 224.560 553.880 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 541.660 224.560 545.200 225.680 ;
  LAYER metal3 ;
  RECT 541.660 224.560 545.200 225.680 ;
  LAYER metal2 ;
  RECT 541.660 224.560 545.200 225.680 ;
  LAYER metal1 ;
  RECT 541.660 224.560 545.200 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 532.980 224.560 536.520 225.680 ;
  LAYER metal3 ;
  RECT 532.980 224.560 536.520 225.680 ;
  LAYER metal2 ;
  RECT 532.980 224.560 536.520 225.680 ;
  LAYER metal1 ;
  RECT 532.980 224.560 536.520 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 489.580 224.560 493.120 225.680 ;
  LAYER metal3 ;
  RECT 489.580 224.560 493.120 225.680 ;
  LAYER metal2 ;
  RECT 489.580 224.560 493.120 225.680 ;
  LAYER metal1 ;
  RECT 489.580 224.560 493.120 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 480.900 224.560 484.440 225.680 ;
  LAYER metal3 ;
  RECT 480.900 224.560 484.440 225.680 ;
  LAYER metal2 ;
  RECT 480.900 224.560 484.440 225.680 ;
  LAYER metal1 ;
  RECT 480.900 224.560 484.440 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 472.220 224.560 475.760 225.680 ;
  LAYER metal3 ;
  RECT 472.220 224.560 475.760 225.680 ;
  LAYER metal2 ;
  RECT 472.220 224.560 475.760 225.680 ;
  LAYER metal1 ;
  RECT 472.220 224.560 475.760 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 463.540 224.560 467.080 225.680 ;
  LAYER metal3 ;
  RECT 463.540 224.560 467.080 225.680 ;
  LAYER metal2 ;
  RECT 463.540 224.560 467.080 225.680 ;
  LAYER metal1 ;
  RECT 463.540 224.560 467.080 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 454.860 224.560 458.400 225.680 ;
  LAYER metal3 ;
  RECT 454.860 224.560 458.400 225.680 ;
  LAYER metal2 ;
  RECT 454.860 224.560 458.400 225.680 ;
  LAYER metal1 ;
  RECT 454.860 224.560 458.400 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 446.180 224.560 449.720 225.680 ;
  LAYER metal3 ;
  RECT 446.180 224.560 449.720 225.680 ;
  LAYER metal2 ;
  RECT 446.180 224.560 449.720 225.680 ;
  LAYER metal1 ;
  RECT 446.180 224.560 449.720 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 402.780 224.560 406.320 225.680 ;
  LAYER metal3 ;
  RECT 402.780 224.560 406.320 225.680 ;
  LAYER metal2 ;
  RECT 402.780 224.560 406.320 225.680 ;
  LAYER metal1 ;
  RECT 402.780 224.560 406.320 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 394.100 224.560 397.640 225.680 ;
  LAYER metal3 ;
  RECT 394.100 224.560 397.640 225.680 ;
  LAYER metal2 ;
  RECT 394.100 224.560 397.640 225.680 ;
  LAYER metal1 ;
  RECT 394.100 224.560 397.640 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 385.420 224.560 388.960 225.680 ;
  LAYER metal3 ;
  RECT 385.420 224.560 388.960 225.680 ;
  LAYER metal2 ;
  RECT 385.420 224.560 388.960 225.680 ;
  LAYER metal1 ;
  RECT 385.420 224.560 388.960 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 376.740 224.560 380.280 225.680 ;
  LAYER metal3 ;
  RECT 376.740 224.560 380.280 225.680 ;
  LAYER metal2 ;
  RECT 376.740 224.560 380.280 225.680 ;
  LAYER metal1 ;
  RECT 376.740 224.560 380.280 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 368.060 224.560 371.600 225.680 ;
  LAYER metal3 ;
  RECT 368.060 224.560 371.600 225.680 ;
  LAYER metal2 ;
  RECT 368.060 224.560 371.600 225.680 ;
  LAYER metal1 ;
  RECT 368.060 224.560 371.600 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 359.380 224.560 362.920 225.680 ;
  LAYER metal3 ;
  RECT 359.380 224.560 362.920 225.680 ;
  LAYER metal2 ;
  RECT 359.380 224.560 362.920 225.680 ;
  LAYER metal1 ;
  RECT 359.380 224.560 362.920 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.980 224.560 319.520 225.680 ;
  LAYER metal3 ;
  RECT 315.980 224.560 319.520 225.680 ;
  LAYER metal2 ;
  RECT 315.980 224.560 319.520 225.680 ;
  LAYER metal1 ;
  RECT 315.980 224.560 319.520 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 307.300 224.560 310.840 225.680 ;
  LAYER metal3 ;
  RECT 307.300 224.560 310.840 225.680 ;
  LAYER metal2 ;
  RECT 307.300 224.560 310.840 225.680 ;
  LAYER metal1 ;
  RECT 307.300 224.560 310.840 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 298.620 224.560 302.160 225.680 ;
  LAYER metal3 ;
  RECT 298.620 224.560 302.160 225.680 ;
  LAYER metal2 ;
  RECT 298.620 224.560 302.160 225.680 ;
  LAYER metal1 ;
  RECT 298.620 224.560 302.160 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 289.940 224.560 293.480 225.680 ;
  LAYER metal3 ;
  RECT 289.940 224.560 293.480 225.680 ;
  LAYER metal2 ;
  RECT 289.940 224.560 293.480 225.680 ;
  LAYER metal1 ;
  RECT 289.940 224.560 293.480 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 281.260 224.560 284.800 225.680 ;
  LAYER metal3 ;
  RECT 281.260 224.560 284.800 225.680 ;
  LAYER metal2 ;
  RECT 281.260 224.560 284.800 225.680 ;
  LAYER metal1 ;
  RECT 281.260 224.560 284.800 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 272.580 224.560 276.120 225.680 ;
  LAYER metal3 ;
  RECT 272.580 224.560 276.120 225.680 ;
  LAYER metal2 ;
  RECT 272.580 224.560 276.120 225.680 ;
  LAYER metal1 ;
  RECT 272.580 224.560 276.120 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 229.180 224.560 232.720 225.680 ;
  LAYER metal3 ;
  RECT 229.180 224.560 232.720 225.680 ;
  LAYER metal2 ;
  RECT 229.180 224.560 232.720 225.680 ;
  LAYER metal1 ;
  RECT 229.180 224.560 232.720 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 220.500 224.560 224.040 225.680 ;
  LAYER metal3 ;
  RECT 220.500 224.560 224.040 225.680 ;
  LAYER metal2 ;
  RECT 220.500 224.560 224.040 225.680 ;
  LAYER metal1 ;
  RECT 220.500 224.560 224.040 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 211.820 224.560 215.360 225.680 ;
  LAYER metal3 ;
  RECT 211.820 224.560 215.360 225.680 ;
  LAYER metal2 ;
  RECT 211.820 224.560 215.360 225.680 ;
  LAYER metal1 ;
  RECT 211.820 224.560 215.360 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 203.140 224.560 206.680 225.680 ;
  LAYER metal3 ;
  RECT 203.140 224.560 206.680 225.680 ;
  LAYER metal2 ;
  RECT 203.140 224.560 206.680 225.680 ;
  LAYER metal1 ;
  RECT 203.140 224.560 206.680 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 194.460 224.560 198.000 225.680 ;
  LAYER metal3 ;
  RECT 194.460 224.560 198.000 225.680 ;
  LAYER metal2 ;
  RECT 194.460 224.560 198.000 225.680 ;
  LAYER metal1 ;
  RECT 194.460 224.560 198.000 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 185.780 224.560 189.320 225.680 ;
  LAYER metal3 ;
  RECT 185.780 224.560 189.320 225.680 ;
  LAYER metal2 ;
  RECT 185.780 224.560 189.320 225.680 ;
  LAYER metal1 ;
  RECT 185.780 224.560 189.320 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 142.380 224.560 145.920 225.680 ;
  LAYER metal3 ;
  RECT 142.380 224.560 145.920 225.680 ;
  LAYER metal2 ;
  RECT 142.380 224.560 145.920 225.680 ;
  LAYER metal1 ;
  RECT 142.380 224.560 145.920 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 133.700 224.560 137.240 225.680 ;
  LAYER metal3 ;
  RECT 133.700 224.560 137.240 225.680 ;
  LAYER metal2 ;
  RECT 133.700 224.560 137.240 225.680 ;
  LAYER metal1 ;
  RECT 133.700 224.560 137.240 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 125.020 224.560 128.560 225.680 ;
  LAYER metal3 ;
  RECT 125.020 224.560 128.560 225.680 ;
  LAYER metal2 ;
  RECT 125.020 224.560 128.560 225.680 ;
  LAYER metal1 ;
  RECT 125.020 224.560 128.560 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 116.340 224.560 119.880 225.680 ;
  LAYER metal3 ;
  RECT 116.340 224.560 119.880 225.680 ;
  LAYER metal2 ;
  RECT 116.340 224.560 119.880 225.680 ;
  LAYER metal1 ;
  RECT 116.340 224.560 119.880 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 107.660 224.560 111.200 225.680 ;
  LAYER metal3 ;
  RECT 107.660 224.560 111.200 225.680 ;
  LAYER metal2 ;
  RECT 107.660 224.560 111.200 225.680 ;
  LAYER metal1 ;
  RECT 107.660 224.560 111.200 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 98.980 224.560 102.520 225.680 ;
  LAYER metal3 ;
  RECT 98.980 224.560 102.520 225.680 ;
  LAYER metal2 ;
  RECT 98.980 224.560 102.520 225.680 ;
  LAYER metal1 ;
  RECT 98.980 224.560 102.520 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 55.580 224.560 59.120 225.680 ;
  LAYER metal3 ;
  RECT 55.580 224.560 59.120 225.680 ;
  LAYER metal2 ;
  RECT 55.580 224.560 59.120 225.680 ;
  LAYER metal1 ;
  RECT 55.580 224.560 59.120 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 46.900 224.560 50.440 225.680 ;
  LAYER metal3 ;
  RECT 46.900 224.560 50.440 225.680 ;
  LAYER metal2 ;
  RECT 46.900 224.560 50.440 225.680 ;
  LAYER metal1 ;
  RECT 46.900 224.560 50.440 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 38.220 224.560 41.760 225.680 ;
  LAYER metal3 ;
  RECT 38.220 224.560 41.760 225.680 ;
  LAYER metal2 ;
  RECT 38.220 224.560 41.760 225.680 ;
  LAYER metal1 ;
  RECT 38.220 224.560 41.760 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 29.540 224.560 33.080 225.680 ;
  LAYER metal3 ;
  RECT 29.540 224.560 33.080 225.680 ;
  LAYER metal2 ;
  RECT 29.540 224.560 33.080 225.680 ;
  LAYER metal1 ;
  RECT 29.540 224.560 33.080 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 20.860 224.560 24.400 225.680 ;
  LAYER metal3 ;
  RECT 20.860 224.560 24.400 225.680 ;
  LAYER metal2 ;
  RECT 20.860 224.560 24.400 225.680 ;
  LAYER metal1 ;
  RECT 20.860 224.560 24.400 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 12.180 224.560 15.720 225.680 ;
  LAYER metal3 ;
  RECT 12.180 224.560 15.720 225.680 ;
  LAYER metal2 ;
  RECT 12.180 224.560 15.720 225.680 ;
  LAYER metal1 ;
  RECT 12.180 224.560 15.720 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 767.960 0.000 771.500 1.120 ;
  LAYER metal3 ;
  RECT 767.960 0.000 771.500 1.120 ;
  LAYER metal2 ;
  RECT 767.960 0.000 771.500 1.120 ;
  LAYER metal1 ;
  RECT 767.960 0.000 771.500 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 746.260 0.000 749.800 1.120 ;
  LAYER metal3 ;
  RECT 746.260 0.000 749.800 1.120 ;
  LAYER metal2 ;
  RECT 746.260 0.000 749.800 1.120 ;
  LAYER metal1 ;
  RECT 746.260 0.000 749.800 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 729.520 0.000 733.060 1.120 ;
  LAYER metal3 ;
  RECT 729.520 0.000 733.060 1.120 ;
  LAYER metal2 ;
  RECT 729.520 0.000 733.060 1.120 ;
  LAYER metal1 ;
  RECT 729.520 0.000 733.060 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 702.860 0.000 706.400 1.120 ;
  LAYER metal3 ;
  RECT 702.860 0.000 706.400 1.120 ;
  LAYER metal2 ;
  RECT 702.860 0.000 706.400 1.120 ;
  LAYER metal1 ;
  RECT 702.860 0.000 706.400 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 681.160 0.000 684.700 1.120 ;
  LAYER metal3 ;
  RECT 681.160 0.000 684.700 1.120 ;
  LAYER metal2 ;
  RECT 681.160 0.000 684.700 1.120 ;
  LAYER metal1 ;
  RECT 681.160 0.000 684.700 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 568.320 0.000 571.860 1.120 ;
  LAYER metal3 ;
  RECT 568.320 0.000 571.860 1.120 ;
  LAYER metal2 ;
  RECT 568.320 0.000 571.860 1.120 ;
  LAYER metal1 ;
  RECT 568.320 0.000 571.860 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 546.620 0.000 550.160 1.120 ;
  LAYER metal3 ;
  RECT 546.620 0.000 550.160 1.120 ;
  LAYER metal2 ;
  RECT 546.620 0.000 550.160 1.120 ;
  LAYER metal1 ;
  RECT 546.620 0.000 550.160 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 519.960 0.000 523.500 1.120 ;
  LAYER metal3 ;
  RECT 519.960 0.000 523.500 1.120 ;
  LAYER metal2 ;
  RECT 519.960 0.000 523.500 1.120 ;
  LAYER metal1 ;
  RECT 519.960 0.000 523.500 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 503.220 0.000 506.760 1.120 ;
  LAYER metal3 ;
  RECT 503.220 0.000 506.760 1.120 ;
  LAYER metal2 ;
  RECT 503.220 0.000 506.760 1.120 ;
  LAYER metal1 ;
  RECT 503.220 0.000 506.760 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 476.560 0.000 480.100 1.120 ;
  LAYER metal3 ;
  RECT 476.560 0.000 480.100 1.120 ;
  LAYER metal2 ;
  RECT 476.560 0.000 480.100 1.120 ;
  LAYER metal1 ;
  RECT 476.560 0.000 480.100 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 454.860 0.000 458.400 1.120 ;
  LAYER metal3 ;
  RECT 454.860 0.000 458.400 1.120 ;
  LAYER metal2 ;
  RECT 454.860 0.000 458.400 1.120 ;
  LAYER metal1 ;
  RECT 454.860 0.000 458.400 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 352.560 0.000 356.100 1.120 ;
  LAYER metal3 ;
  RECT 352.560 0.000 356.100 1.120 ;
  LAYER metal2 ;
  RECT 352.560 0.000 356.100 1.120 ;
  LAYER metal1 ;
  RECT 352.560 0.000 356.100 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 339.540 0.000 343.080 1.120 ;
  LAYER metal3 ;
  RECT 339.540 0.000 343.080 1.120 ;
  LAYER metal2 ;
  RECT 339.540 0.000 343.080 1.120 ;
  LAYER metal1 ;
  RECT 339.540 0.000 343.080 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 318.460 0.000 322.000 1.120 ;
  LAYER metal3 ;
  RECT 318.460 0.000 322.000 1.120 ;
  LAYER metal2 ;
  RECT 318.460 0.000 322.000 1.120 ;
  LAYER metal1 ;
  RECT 318.460 0.000 322.000 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 296.760 0.000 300.300 1.120 ;
  LAYER metal3 ;
  RECT 296.760 0.000 300.300 1.120 ;
  LAYER metal2 ;
  RECT 296.760 0.000 300.300 1.120 ;
  LAYER metal1 ;
  RECT 296.760 0.000 300.300 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 270.100 0.000 273.640 1.120 ;
  LAYER metal3 ;
  RECT 270.100 0.000 273.640 1.120 ;
  LAYER metal2 ;
  RECT 270.100 0.000 273.640 1.120 ;
  LAYER metal1 ;
  RECT 270.100 0.000 273.640 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER metal3 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER metal2 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER metal1 ;
  RECT 253.360 0.000 256.900 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER metal3 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER metal2 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER metal1 ;
  RECT 139.900 0.000 143.440 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER metal3 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER metal2 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER metal1 ;
  RECT 113.860 0.000 117.400 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER metal3 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER metal2 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER metal1 ;
  RECT 92.160 0.000 95.700 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal3 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal2 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal1 ;
  RECT 70.460 0.000 74.000 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER metal3 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER metal2 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER metal1 ;
  RECT 43.800 0.000 47.340 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal3 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal2 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal1 ;
  RECT 27.060 0.000 30.600 1.120 ;
 END
END GND
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal4 ;
  RECT 777.600 204.180 778.720 207.420 ;
  LAYER metal3 ;
  RECT 777.600 204.180 778.720 207.420 ;
  LAYER metal2 ;
  RECT 777.600 204.180 778.720 207.420 ;
  LAYER metal1 ;
  RECT 777.600 204.180 778.720 207.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 196.340 778.720 199.580 ;
  LAYER metal3 ;
  RECT 777.600 196.340 778.720 199.580 ;
  LAYER metal2 ;
  RECT 777.600 196.340 778.720 199.580 ;
  LAYER metal1 ;
  RECT 777.600 196.340 778.720 199.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 188.500 778.720 191.740 ;
  LAYER metal3 ;
  RECT 777.600 188.500 778.720 191.740 ;
  LAYER metal2 ;
  RECT 777.600 188.500 778.720 191.740 ;
  LAYER metal1 ;
  RECT 777.600 188.500 778.720 191.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 180.660 778.720 183.900 ;
  LAYER metal3 ;
  RECT 777.600 180.660 778.720 183.900 ;
  LAYER metal2 ;
  RECT 777.600 180.660 778.720 183.900 ;
  LAYER metal1 ;
  RECT 777.600 180.660 778.720 183.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 172.820 778.720 176.060 ;
  LAYER metal3 ;
  RECT 777.600 172.820 778.720 176.060 ;
  LAYER metal2 ;
  RECT 777.600 172.820 778.720 176.060 ;
  LAYER metal1 ;
  RECT 777.600 172.820 778.720 176.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 164.980 778.720 168.220 ;
  LAYER metal3 ;
  RECT 777.600 164.980 778.720 168.220 ;
  LAYER metal2 ;
  RECT 777.600 164.980 778.720 168.220 ;
  LAYER metal1 ;
  RECT 777.600 164.980 778.720 168.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 125.780 778.720 129.020 ;
  LAYER metal3 ;
  RECT 777.600 125.780 778.720 129.020 ;
  LAYER metal2 ;
  RECT 777.600 125.780 778.720 129.020 ;
  LAYER metal1 ;
  RECT 777.600 125.780 778.720 129.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 117.940 778.720 121.180 ;
  LAYER metal3 ;
  RECT 777.600 117.940 778.720 121.180 ;
  LAYER metal2 ;
  RECT 777.600 117.940 778.720 121.180 ;
  LAYER metal1 ;
  RECT 777.600 117.940 778.720 121.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 110.100 778.720 113.340 ;
  LAYER metal3 ;
  RECT 777.600 110.100 778.720 113.340 ;
  LAYER metal2 ;
  RECT 777.600 110.100 778.720 113.340 ;
  LAYER metal1 ;
  RECT 777.600 110.100 778.720 113.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 102.260 778.720 105.500 ;
  LAYER metal3 ;
  RECT 777.600 102.260 778.720 105.500 ;
  LAYER metal2 ;
  RECT 777.600 102.260 778.720 105.500 ;
  LAYER metal1 ;
  RECT 777.600 102.260 778.720 105.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 94.420 778.720 97.660 ;
  LAYER metal3 ;
  RECT 777.600 94.420 778.720 97.660 ;
  LAYER metal2 ;
  RECT 777.600 94.420 778.720 97.660 ;
  LAYER metal1 ;
  RECT 777.600 94.420 778.720 97.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 86.580 778.720 89.820 ;
  LAYER metal3 ;
  RECT 777.600 86.580 778.720 89.820 ;
  LAYER metal2 ;
  RECT 777.600 86.580 778.720 89.820 ;
  LAYER metal1 ;
  RECT 777.600 86.580 778.720 89.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 47.380 778.720 50.620 ;
  LAYER metal3 ;
  RECT 777.600 47.380 778.720 50.620 ;
  LAYER metal2 ;
  RECT 777.600 47.380 778.720 50.620 ;
  LAYER metal1 ;
  RECT 777.600 47.380 778.720 50.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 39.540 778.720 42.780 ;
  LAYER metal3 ;
  RECT 777.600 39.540 778.720 42.780 ;
  LAYER metal2 ;
  RECT 777.600 39.540 778.720 42.780 ;
  LAYER metal1 ;
  RECT 777.600 39.540 778.720 42.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 31.700 778.720 34.940 ;
  LAYER metal3 ;
  RECT 777.600 31.700 778.720 34.940 ;
  LAYER metal2 ;
  RECT 777.600 31.700 778.720 34.940 ;
  LAYER metal1 ;
  RECT 777.600 31.700 778.720 34.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 23.860 778.720 27.100 ;
  LAYER metal3 ;
  RECT 777.600 23.860 778.720 27.100 ;
  LAYER metal2 ;
  RECT 777.600 23.860 778.720 27.100 ;
  LAYER metal1 ;
  RECT 777.600 23.860 778.720 27.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 16.020 778.720 19.260 ;
  LAYER metal3 ;
  RECT 777.600 16.020 778.720 19.260 ;
  LAYER metal2 ;
  RECT 777.600 16.020 778.720 19.260 ;
  LAYER metal1 ;
  RECT 777.600 16.020 778.720 19.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 777.600 8.180 778.720 11.420 ;
  LAYER metal3 ;
  RECT 777.600 8.180 778.720 11.420 ;
  LAYER metal2 ;
  RECT 777.600 8.180 778.720 11.420 ;
  LAYER metal1 ;
  RECT 777.600 8.180 778.720 11.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER metal3 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER metal2 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER metal1 ;
  RECT 0.000 204.180 1.120 207.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER metal3 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER metal2 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER metal1 ;
  RECT 0.000 196.340 1.120 199.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER metal3 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER metal2 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER metal1 ;
  RECT 0.000 188.500 1.120 191.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER metal3 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER metal2 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER metal1 ;
  RECT 0.000 180.660 1.120 183.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER metal3 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER metal2 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER metal1 ;
  RECT 0.000 172.820 1.120 176.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER metal3 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER metal2 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER metal1 ;
  RECT 0.000 164.980 1.120 168.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal3 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal2 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal1 ;
  RECT 0.000 125.780 1.120 129.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal3 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal2 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal1 ;
  RECT 0.000 117.940 1.120 121.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal3 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal2 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal1 ;
  RECT 0.000 110.100 1.120 113.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal3 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal2 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal1 ;
  RECT 0.000 102.260 1.120 105.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal3 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal2 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal1 ;
  RECT 0.000 94.420 1.120 97.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal3 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal2 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal1 ;
  RECT 0.000 86.580 1.120 89.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal3 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal2 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal1 ;
  RECT 0.000 47.380 1.120 50.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal3 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal2 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal1 ;
  RECT 0.000 39.540 1.120 42.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal3 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal2 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal1 ;
  RECT 0.000 31.700 1.120 34.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal3 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal2 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal1 ;
  RECT 0.000 23.860 1.120 27.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal3 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal2 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal1 ;
  RECT 0.000 16.020 1.120 19.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal3 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal2 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal1 ;
  RECT 0.000 8.180 1.120 11.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 745.640 224.560 749.180 225.680 ;
  LAYER metal3 ;
  RECT 745.640 224.560 749.180 225.680 ;
  LAYER metal2 ;
  RECT 745.640 224.560 749.180 225.680 ;
  LAYER metal1 ;
  RECT 745.640 224.560 749.180 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 736.960 224.560 740.500 225.680 ;
  LAYER metal3 ;
  RECT 736.960 224.560 740.500 225.680 ;
  LAYER metal2 ;
  RECT 736.960 224.560 740.500 225.680 ;
  LAYER metal1 ;
  RECT 736.960 224.560 740.500 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 728.280 224.560 731.820 225.680 ;
  LAYER metal3 ;
  RECT 728.280 224.560 731.820 225.680 ;
  LAYER metal2 ;
  RECT 728.280 224.560 731.820 225.680 ;
  LAYER metal1 ;
  RECT 728.280 224.560 731.820 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 719.600 224.560 723.140 225.680 ;
  LAYER metal3 ;
  RECT 719.600 224.560 723.140 225.680 ;
  LAYER metal2 ;
  RECT 719.600 224.560 723.140 225.680 ;
  LAYER metal1 ;
  RECT 719.600 224.560 723.140 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 710.920 224.560 714.460 225.680 ;
  LAYER metal3 ;
  RECT 710.920 224.560 714.460 225.680 ;
  LAYER metal2 ;
  RECT 710.920 224.560 714.460 225.680 ;
  LAYER metal1 ;
  RECT 710.920 224.560 714.460 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 702.240 224.560 705.780 225.680 ;
  LAYER metal3 ;
  RECT 702.240 224.560 705.780 225.680 ;
  LAYER metal2 ;
  RECT 702.240 224.560 705.780 225.680 ;
  LAYER metal1 ;
  RECT 702.240 224.560 705.780 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 658.840 224.560 662.380 225.680 ;
  LAYER metal3 ;
  RECT 658.840 224.560 662.380 225.680 ;
  LAYER metal2 ;
  RECT 658.840 224.560 662.380 225.680 ;
  LAYER metal1 ;
  RECT 658.840 224.560 662.380 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 650.160 224.560 653.700 225.680 ;
  LAYER metal3 ;
  RECT 650.160 224.560 653.700 225.680 ;
  LAYER metal2 ;
  RECT 650.160 224.560 653.700 225.680 ;
  LAYER metal1 ;
  RECT 650.160 224.560 653.700 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 641.480 224.560 645.020 225.680 ;
  LAYER metal3 ;
  RECT 641.480 224.560 645.020 225.680 ;
  LAYER metal2 ;
  RECT 641.480 224.560 645.020 225.680 ;
  LAYER metal1 ;
  RECT 641.480 224.560 645.020 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 632.800 224.560 636.340 225.680 ;
  LAYER metal3 ;
  RECT 632.800 224.560 636.340 225.680 ;
  LAYER metal2 ;
  RECT 632.800 224.560 636.340 225.680 ;
  LAYER metal1 ;
  RECT 632.800 224.560 636.340 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 624.120 224.560 627.660 225.680 ;
  LAYER metal3 ;
  RECT 624.120 224.560 627.660 225.680 ;
  LAYER metal2 ;
  RECT 624.120 224.560 627.660 225.680 ;
  LAYER metal1 ;
  RECT 624.120 224.560 627.660 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 615.440 224.560 618.980 225.680 ;
  LAYER metal3 ;
  RECT 615.440 224.560 618.980 225.680 ;
  LAYER metal2 ;
  RECT 615.440 224.560 618.980 225.680 ;
  LAYER metal1 ;
  RECT 615.440 224.560 618.980 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 572.040 224.560 575.580 225.680 ;
  LAYER metal3 ;
  RECT 572.040 224.560 575.580 225.680 ;
  LAYER metal2 ;
  RECT 572.040 224.560 575.580 225.680 ;
  LAYER metal1 ;
  RECT 572.040 224.560 575.580 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 563.360 224.560 566.900 225.680 ;
  LAYER metal3 ;
  RECT 563.360 224.560 566.900 225.680 ;
  LAYER metal2 ;
  RECT 563.360 224.560 566.900 225.680 ;
  LAYER metal1 ;
  RECT 563.360 224.560 566.900 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 554.680 224.560 558.220 225.680 ;
  LAYER metal3 ;
  RECT 554.680 224.560 558.220 225.680 ;
  LAYER metal2 ;
  RECT 554.680 224.560 558.220 225.680 ;
  LAYER metal1 ;
  RECT 554.680 224.560 558.220 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 546.000 224.560 549.540 225.680 ;
  LAYER metal3 ;
  RECT 546.000 224.560 549.540 225.680 ;
  LAYER metal2 ;
  RECT 546.000 224.560 549.540 225.680 ;
  LAYER metal1 ;
  RECT 546.000 224.560 549.540 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 537.320 224.560 540.860 225.680 ;
  LAYER metal3 ;
  RECT 537.320 224.560 540.860 225.680 ;
  LAYER metal2 ;
  RECT 537.320 224.560 540.860 225.680 ;
  LAYER metal1 ;
  RECT 537.320 224.560 540.860 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 528.640 224.560 532.180 225.680 ;
  LAYER metal3 ;
  RECT 528.640 224.560 532.180 225.680 ;
  LAYER metal2 ;
  RECT 528.640 224.560 532.180 225.680 ;
  LAYER metal1 ;
  RECT 528.640 224.560 532.180 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 485.240 224.560 488.780 225.680 ;
  LAYER metal3 ;
  RECT 485.240 224.560 488.780 225.680 ;
  LAYER metal2 ;
  RECT 485.240 224.560 488.780 225.680 ;
  LAYER metal1 ;
  RECT 485.240 224.560 488.780 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 476.560 224.560 480.100 225.680 ;
  LAYER metal3 ;
  RECT 476.560 224.560 480.100 225.680 ;
  LAYER metal2 ;
  RECT 476.560 224.560 480.100 225.680 ;
  LAYER metal1 ;
  RECT 476.560 224.560 480.100 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 467.880 224.560 471.420 225.680 ;
  LAYER metal3 ;
  RECT 467.880 224.560 471.420 225.680 ;
  LAYER metal2 ;
  RECT 467.880 224.560 471.420 225.680 ;
  LAYER metal1 ;
  RECT 467.880 224.560 471.420 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 459.200 224.560 462.740 225.680 ;
  LAYER metal3 ;
  RECT 459.200 224.560 462.740 225.680 ;
  LAYER metal2 ;
  RECT 459.200 224.560 462.740 225.680 ;
  LAYER metal1 ;
  RECT 459.200 224.560 462.740 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 450.520 224.560 454.060 225.680 ;
  LAYER metal3 ;
  RECT 450.520 224.560 454.060 225.680 ;
  LAYER metal2 ;
  RECT 450.520 224.560 454.060 225.680 ;
  LAYER metal1 ;
  RECT 450.520 224.560 454.060 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 441.840 224.560 445.380 225.680 ;
  LAYER metal3 ;
  RECT 441.840 224.560 445.380 225.680 ;
  LAYER metal2 ;
  RECT 441.840 224.560 445.380 225.680 ;
  LAYER metal1 ;
  RECT 441.840 224.560 445.380 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 398.440 224.560 401.980 225.680 ;
  LAYER metal3 ;
  RECT 398.440 224.560 401.980 225.680 ;
  LAYER metal2 ;
  RECT 398.440 224.560 401.980 225.680 ;
  LAYER metal1 ;
  RECT 398.440 224.560 401.980 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 389.760 224.560 393.300 225.680 ;
  LAYER metal3 ;
  RECT 389.760 224.560 393.300 225.680 ;
  LAYER metal2 ;
  RECT 389.760 224.560 393.300 225.680 ;
  LAYER metal1 ;
  RECT 389.760 224.560 393.300 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 381.080 224.560 384.620 225.680 ;
  LAYER metal3 ;
  RECT 381.080 224.560 384.620 225.680 ;
  LAYER metal2 ;
  RECT 381.080 224.560 384.620 225.680 ;
  LAYER metal1 ;
  RECT 381.080 224.560 384.620 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 372.400 224.560 375.940 225.680 ;
  LAYER metal3 ;
  RECT 372.400 224.560 375.940 225.680 ;
  LAYER metal2 ;
  RECT 372.400 224.560 375.940 225.680 ;
  LAYER metal1 ;
  RECT 372.400 224.560 375.940 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 363.720 224.560 367.260 225.680 ;
  LAYER metal3 ;
  RECT 363.720 224.560 367.260 225.680 ;
  LAYER metal2 ;
  RECT 363.720 224.560 367.260 225.680 ;
  LAYER metal1 ;
  RECT 363.720 224.560 367.260 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 355.040 224.560 358.580 225.680 ;
  LAYER metal3 ;
  RECT 355.040 224.560 358.580 225.680 ;
  LAYER metal2 ;
  RECT 355.040 224.560 358.580 225.680 ;
  LAYER metal1 ;
  RECT 355.040 224.560 358.580 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 311.640 224.560 315.180 225.680 ;
  LAYER metal3 ;
  RECT 311.640 224.560 315.180 225.680 ;
  LAYER metal2 ;
  RECT 311.640 224.560 315.180 225.680 ;
  LAYER metal1 ;
  RECT 311.640 224.560 315.180 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 302.960 224.560 306.500 225.680 ;
  LAYER metal3 ;
  RECT 302.960 224.560 306.500 225.680 ;
  LAYER metal2 ;
  RECT 302.960 224.560 306.500 225.680 ;
  LAYER metal1 ;
  RECT 302.960 224.560 306.500 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 294.280 224.560 297.820 225.680 ;
  LAYER metal3 ;
  RECT 294.280 224.560 297.820 225.680 ;
  LAYER metal2 ;
  RECT 294.280 224.560 297.820 225.680 ;
  LAYER metal1 ;
  RECT 294.280 224.560 297.820 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 285.600 224.560 289.140 225.680 ;
  LAYER metal3 ;
  RECT 285.600 224.560 289.140 225.680 ;
  LAYER metal2 ;
  RECT 285.600 224.560 289.140 225.680 ;
  LAYER metal1 ;
  RECT 285.600 224.560 289.140 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 276.920 224.560 280.460 225.680 ;
  LAYER metal3 ;
  RECT 276.920 224.560 280.460 225.680 ;
  LAYER metal2 ;
  RECT 276.920 224.560 280.460 225.680 ;
  LAYER metal1 ;
  RECT 276.920 224.560 280.460 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 268.240 224.560 271.780 225.680 ;
  LAYER metal3 ;
  RECT 268.240 224.560 271.780 225.680 ;
  LAYER metal2 ;
  RECT 268.240 224.560 271.780 225.680 ;
  LAYER metal1 ;
  RECT 268.240 224.560 271.780 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 224.840 224.560 228.380 225.680 ;
  LAYER metal3 ;
  RECT 224.840 224.560 228.380 225.680 ;
  LAYER metal2 ;
  RECT 224.840 224.560 228.380 225.680 ;
  LAYER metal1 ;
  RECT 224.840 224.560 228.380 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 216.160 224.560 219.700 225.680 ;
  LAYER metal3 ;
  RECT 216.160 224.560 219.700 225.680 ;
  LAYER metal2 ;
  RECT 216.160 224.560 219.700 225.680 ;
  LAYER metal1 ;
  RECT 216.160 224.560 219.700 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 207.480 224.560 211.020 225.680 ;
  LAYER metal3 ;
  RECT 207.480 224.560 211.020 225.680 ;
  LAYER metal2 ;
  RECT 207.480 224.560 211.020 225.680 ;
  LAYER metal1 ;
  RECT 207.480 224.560 211.020 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 198.800 224.560 202.340 225.680 ;
  LAYER metal3 ;
  RECT 198.800 224.560 202.340 225.680 ;
  LAYER metal2 ;
  RECT 198.800 224.560 202.340 225.680 ;
  LAYER metal1 ;
  RECT 198.800 224.560 202.340 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 190.120 224.560 193.660 225.680 ;
  LAYER metal3 ;
  RECT 190.120 224.560 193.660 225.680 ;
  LAYER metal2 ;
  RECT 190.120 224.560 193.660 225.680 ;
  LAYER metal1 ;
  RECT 190.120 224.560 193.660 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 181.440 224.560 184.980 225.680 ;
  LAYER metal3 ;
  RECT 181.440 224.560 184.980 225.680 ;
  LAYER metal2 ;
  RECT 181.440 224.560 184.980 225.680 ;
  LAYER metal1 ;
  RECT 181.440 224.560 184.980 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 138.040 224.560 141.580 225.680 ;
  LAYER metal3 ;
  RECT 138.040 224.560 141.580 225.680 ;
  LAYER metal2 ;
  RECT 138.040 224.560 141.580 225.680 ;
  LAYER metal1 ;
  RECT 138.040 224.560 141.580 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 129.360 224.560 132.900 225.680 ;
  LAYER metal3 ;
  RECT 129.360 224.560 132.900 225.680 ;
  LAYER metal2 ;
  RECT 129.360 224.560 132.900 225.680 ;
  LAYER metal1 ;
  RECT 129.360 224.560 132.900 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 120.680 224.560 124.220 225.680 ;
  LAYER metal3 ;
  RECT 120.680 224.560 124.220 225.680 ;
  LAYER metal2 ;
  RECT 120.680 224.560 124.220 225.680 ;
  LAYER metal1 ;
  RECT 120.680 224.560 124.220 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 112.000 224.560 115.540 225.680 ;
  LAYER metal3 ;
  RECT 112.000 224.560 115.540 225.680 ;
  LAYER metal2 ;
  RECT 112.000 224.560 115.540 225.680 ;
  LAYER metal1 ;
  RECT 112.000 224.560 115.540 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 103.320 224.560 106.860 225.680 ;
  LAYER metal3 ;
  RECT 103.320 224.560 106.860 225.680 ;
  LAYER metal2 ;
  RECT 103.320 224.560 106.860 225.680 ;
  LAYER metal1 ;
  RECT 103.320 224.560 106.860 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 94.640 224.560 98.180 225.680 ;
  LAYER metal3 ;
  RECT 94.640 224.560 98.180 225.680 ;
  LAYER metal2 ;
  RECT 94.640 224.560 98.180 225.680 ;
  LAYER metal1 ;
  RECT 94.640 224.560 98.180 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 51.240 224.560 54.780 225.680 ;
  LAYER metal3 ;
  RECT 51.240 224.560 54.780 225.680 ;
  LAYER metal2 ;
  RECT 51.240 224.560 54.780 225.680 ;
  LAYER metal1 ;
  RECT 51.240 224.560 54.780 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 42.560 224.560 46.100 225.680 ;
  LAYER metal3 ;
  RECT 42.560 224.560 46.100 225.680 ;
  LAYER metal2 ;
  RECT 42.560 224.560 46.100 225.680 ;
  LAYER metal1 ;
  RECT 42.560 224.560 46.100 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 33.880 224.560 37.420 225.680 ;
  LAYER metal3 ;
  RECT 33.880 224.560 37.420 225.680 ;
  LAYER metal2 ;
  RECT 33.880 224.560 37.420 225.680 ;
  LAYER metal1 ;
  RECT 33.880 224.560 37.420 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 25.200 224.560 28.740 225.680 ;
  LAYER metal3 ;
  RECT 25.200 224.560 28.740 225.680 ;
  LAYER metal2 ;
  RECT 25.200 224.560 28.740 225.680 ;
  LAYER metal1 ;
  RECT 25.200 224.560 28.740 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 16.520 224.560 20.060 225.680 ;
  LAYER metal3 ;
  RECT 16.520 224.560 20.060 225.680 ;
  LAYER metal2 ;
  RECT 16.520 224.560 20.060 225.680 ;
  LAYER metal1 ;
  RECT 16.520 224.560 20.060 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 7.840 224.560 11.380 225.680 ;
  LAYER metal3 ;
  RECT 7.840 224.560 11.380 225.680 ;
  LAYER metal2 ;
  RECT 7.840 224.560 11.380 225.680 ;
  LAYER metal1 ;
  RECT 7.840 224.560 11.380 225.680 ;
 END
 PORT
  LAYER metal4 ;
  RECT 759.280 0.000 762.820 1.120 ;
  LAYER metal3 ;
  RECT 759.280 0.000 762.820 1.120 ;
  LAYER metal2 ;
  RECT 759.280 0.000 762.820 1.120 ;
  LAYER metal1 ;
  RECT 759.280 0.000 762.820 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 737.580 0.000 741.120 1.120 ;
  LAYER metal3 ;
  RECT 737.580 0.000 741.120 1.120 ;
  LAYER metal2 ;
  RECT 737.580 0.000 741.120 1.120 ;
  LAYER metal1 ;
  RECT 737.580 0.000 741.120 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 715.880 0.000 719.420 1.120 ;
  LAYER metal3 ;
  RECT 715.880 0.000 719.420 1.120 ;
  LAYER metal2 ;
  RECT 715.880 0.000 719.420 1.120 ;
  LAYER metal1 ;
  RECT 715.880 0.000 719.420 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 689.220 0.000 692.760 1.120 ;
  LAYER metal3 ;
  RECT 689.220 0.000 692.760 1.120 ;
  LAYER metal2 ;
  RECT 689.220 0.000 692.760 1.120 ;
  LAYER metal1 ;
  RECT 689.220 0.000 692.760 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 673.100 0.000 676.640 1.120 ;
  LAYER metal3 ;
  RECT 673.100 0.000 676.640 1.120 ;
  LAYER metal2 ;
  RECT 673.100 0.000 676.640 1.120 ;
  LAYER metal1 ;
  RECT 673.100 0.000 676.640 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 559.640 0.000 563.180 1.120 ;
  LAYER metal3 ;
  RECT 559.640 0.000 563.180 1.120 ;
  LAYER metal2 ;
  RECT 559.640 0.000 563.180 1.120 ;
  LAYER metal1 ;
  RECT 559.640 0.000 563.180 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 532.980 0.000 536.520 1.120 ;
  LAYER metal3 ;
  RECT 532.980 0.000 536.520 1.120 ;
  LAYER metal2 ;
  RECT 532.980 0.000 536.520 1.120 ;
  LAYER metal1 ;
  RECT 532.980 0.000 536.520 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 511.900 0.000 515.440 1.120 ;
  LAYER metal3 ;
  RECT 511.900 0.000 515.440 1.120 ;
  LAYER metal2 ;
  RECT 511.900 0.000 515.440 1.120 ;
  LAYER metal1 ;
  RECT 511.900 0.000 515.440 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 490.200 0.000 493.740 1.120 ;
  LAYER metal3 ;
  RECT 490.200 0.000 493.740 1.120 ;
  LAYER metal2 ;
  RECT 490.200 0.000 493.740 1.120 ;
  LAYER metal1 ;
  RECT 490.200 0.000 493.740 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 463.540 0.000 467.080 1.120 ;
  LAYER metal3 ;
  RECT 463.540 0.000 467.080 1.120 ;
  LAYER metal2 ;
  RECT 463.540 0.000 467.080 1.120 ;
  LAYER metal1 ;
  RECT 463.540 0.000 467.080 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 446.800 0.000 450.340 1.120 ;
  LAYER metal3 ;
  RECT 446.800 0.000 450.340 1.120 ;
  LAYER metal2 ;
  RECT 446.800 0.000 450.340 1.120 ;
  LAYER metal1 ;
  RECT 446.800 0.000 450.340 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 348.220 0.000 351.760 1.120 ;
  LAYER metal3 ;
  RECT 348.220 0.000 351.760 1.120 ;
  LAYER metal2 ;
  RECT 348.220 0.000 351.760 1.120 ;
  LAYER metal1 ;
  RECT 348.220 0.000 351.760 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 326.520 0.000 330.060 1.120 ;
  LAYER metal3 ;
  RECT 326.520 0.000 330.060 1.120 ;
  LAYER metal2 ;
  RECT 326.520 0.000 330.060 1.120 ;
  LAYER metal1 ;
  RECT 326.520 0.000 330.060 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 309.780 0.000 313.320 1.120 ;
  LAYER metal3 ;
  RECT 309.780 0.000 313.320 1.120 ;
  LAYER metal2 ;
  RECT 309.780 0.000 313.320 1.120 ;
  LAYER metal1 ;
  RECT 309.780 0.000 313.320 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER metal3 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER metal2 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER metal1 ;
  RECT 283.120 0.000 286.660 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER metal3 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER metal2 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER metal1 ;
  RECT 261.420 0.000 264.960 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER metal3 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER metal2 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER metal1 ;
  RECT 239.720 0.000 243.260 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER metal3 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER metal2 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER metal1 ;
  RECT 126.880 0.000 130.420 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER metal3 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER metal2 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER metal1 ;
  RECT 100.220 0.000 103.760 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER metal3 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER metal2 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER metal1 ;
  RECT 83.480 0.000 87.020 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER metal3 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER metal2 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER metal1 ;
  RECT 56.820 0.000 60.360 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal3 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal2 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal1 ;
  RECT 35.740 0.000 39.280 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal3 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal2 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal1 ;
  RECT 14.040 0.000 17.580 1.120 ;
 END
END VCC
PIN DO47
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 765.760 0.000 766.880 1.120 ;
  LAYER metal3 ;
  RECT 765.760 0.000 766.880 1.120 ;
  LAYER metal2 ;
  RECT 765.760 0.000 766.880 1.120 ;
  LAYER metal1 ;
  RECT 765.760 0.000 766.880 1.120 ;
 END
END DO47
PIN DI47
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 757.080 0.000 758.200 1.120 ;
  LAYER metal3 ;
  RECT 757.080 0.000 758.200 1.120 ;
  LAYER metal2 ;
  RECT 757.080 0.000 758.200 1.120 ;
  LAYER metal1 ;
  RECT 757.080 0.000 758.200 1.120 ;
 END
END DI47
PIN DO46
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 752.120 0.000 753.240 1.120 ;
  LAYER metal3 ;
  RECT 752.120 0.000 753.240 1.120 ;
  LAYER metal2 ;
  RECT 752.120 0.000 753.240 1.120 ;
  LAYER metal1 ;
  RECT 752.120 0.000 753.240 1.120 ;
 END
END DO46
PIN DI46
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 744.060 0.000 745.180 1.120 ;
  LAYER metal3 ;
  RECT 744.060 0.000 745.180 1.120 ;
  LAYER metal2 ;
  RECT 744.060 0.000 745.180 1.120 ;
  LAYER metal1 ;
  RECT 744.060 0.000 745.180 1.120 ;
 END
END DI46
PIN DO45
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 735.380 0.000 736.500 1.120 ;
  LAYER metal3 ;
  RECT 735.380 0.000 736.500 1.120 ;
  LAYER metal2 ;
  RECT 735.380 0.000 736.500 1.120 ;
  LAYER metal1 ;
  RECT 735.380 0.000 736.500 1.120 ;
 END
END DO45
PIN DI45
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 727.320 0.000 728.440 1.120 ;
  LAYER metal3 ;
  RECT 727.320 0.000 728.440 1.120 ;
  LAYER metal2 ;
  RECT 727.320 0.000 728.440 1.120 ;
  LAYER metal1 ;
  RECT 727.320 0.000 728.440 1.120 ;
 END
END DI45
PIN DO44
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 722.360 0.000 723.480 1.120 ;
  LAYER metal3 ;
  RECT 722.360 0.000 723.480 1.120 ;
  LAYER metal2 ;
  RECT 722.360 0.000 723.480 1.120 ;
  LAYER metal1 ;
  RECT 722.360 0.000 723.480 1.120 ;
 END
END DO44
PIN DI44
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 713.680 0.000 714.800 1.120 ;
  LAYER metal3 ;
  RECT 713.680 0.000 714.800 1.120 ;
  LAYER metal2 ;
  RECT 713.680 0.000 714.800 1.120 ;
  LAYER metal1 ;
  RECT 713.680 0.000 714.800 1.120 ;
 END
END DI44
PIN DO43
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 708.720 0.000 709.840 1.120 ;
  LAYER metal3 ;
  RECT 708.720 0.000 709.840 1.120 ;
  LAYER metal2 ;
  RECT 708.720 0.000 709.840 1.120 ;
  LAYER metal1 ;
  RECT 708.720 0.000 709.840 1.120 ;
 END
END DO43
PIN DI43
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 700.660 0.000 701.780 1.120 ;
  LAYER metal3 ;
  RECT 700.660 0.000 701.780 1.120 ;
  LAYER metal2 ;
  RECT 700.660 0.000 701.780 1.120 ;
  LAYER metal1 ;
  RECT 700.660 0.000 701.780 1.120 ;
 END
END DI43
PIN DO42
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 695.700 0.000 696.820 1.120 ;
  LAYER metal3 ;
  RECT 695.700 0.000 696.820 1.120 ;
  LAYER metal2 ;
  RECT 695.700 0.000 696.820 1.120 ;
  LAYER metal1 ;
  RECT 695.700 0.000 696.820 1.120 ;
 END
END DO42
PIN DI42
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 687.020 0.000 688.140 1.120 ;
  LAYER metal3 ;
  RECT 687.020 0.000 688.140 1.120 ;
  LAYER metal2 ;
  RECT 687.020 0.000 688.140 1.120 ;
  LAYER metal1 ;
  RECT 687.020 0.000 688.140 1.120 ;
 END
END DI42
PIN DO41
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 678.960 0.000 680.080 1.120 ;
  LAYER metal3 ;
  RECT 678.960 0.000 680.080 1.120 ;
  LAYER metal2 ;
  RECT 678.960 0.000 680.080 1.120 ;
  LAYER metal1 ;
  RECT 678.960 0.000 680.080 1.120 ;
 END
END DO41
PIN DI41
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 670.900 0.000 672.020 1.120 ;
  LAYER metal3 ;
  RECT 670.900 0.000 672.020 1.120 ;
  LAYER metal2 ;
  RECT 670.900 0.000 672.020 1.120 ;
  LAYER metal1 ;
  RECT 670.900 0.000 672.020 1.120 ;
 END
END DI41
PIN DO40
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 665.940 0.000 667.060 1.120 ;
  LAYER metal3 ;
  RECT 665.940 0.000 667.060 1.120 ;
  LAYER metal2 ;
  RECT 665.940 0.000 667.060 1.120 ;
  LAYER metal1 ;
  RECT 665.940 0.000 667.060 1.120 ;
 END
END DO40
PIN DI40
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 657.260 0.000 658.380 1.120 ;
  LAYER metal3 ;
  RECT 657.260 0.000 658.380 1.120 ;
  LAYER metal2 ;
  RECT 657.260 0.000 658.380 1.120 ;
  LAYER metal1 ;
  RECT 657.260 0.000 658.380 1.120 ;
 END
END DI40
PIN DO39
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 652.300 0.000 653.420 1.120 ;
  LAYER metal3 ;
  RECT 652.300 0.000 653.420 1.120 ;
  LAYER metal2 ;
  RECT 652.300 0.000 653.420 1.120 ;
  LAYER metal1 ;
  RECT 652.300 0.000 653.420 1.120 ;
 END
END DO39
PIN DI39
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 644.240 0.000 645.360 1.120 ;
  LAYER metal3 ;
  RECT 644.240 0.000 645.360 1.120 ;
  LAYER metal2 ;
  RECT 644.240 0.000 645.360 1.120 ;
  LAYER metal1 ;
  RECT 644.240 0.000 645.360 1.120 ;
 END
END DI39
PIN DO38
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 639.280 0.000 640.400 1.120 ;
  LAYER metal3 ;
  RECT 639.280 0.000 640.400 1.120 ;
  LAYER metal2 ;
  RECT 639.280 0.000 640.400 1.120 ;
  LAYER metal1 ;
  RECT 639.280 0.000 640.400 1.120 ;
 END
END DO38
PIN DI38
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 630.600 0.000 631.720 1.120 ;
  LAYER metal3 ;
  RECT 630.600 0.000 631.720 1.120 ;
  LAYER metal2 ;
  RECT 630.600 0.000 631.720 1.120 ;
  LAYER metal1 ;
  RECT 630.600 0.000 631.720 1.120 ;
 END
END DI38
PIN DO37
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 622.540 0.000 623.660 1.120 ;
  LAYER metal3 ;
  RECT 622.540 0.000 623.660 1.120 ;
  LAYER metal2 ;
  RECT 622.540 0.000 623.660 1.120 ;
  LAYER metal1 ;
  RECT 622.540 0.000 623.660 1.120 ;
 END
END DO37
PIN DI37
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 613.860 0.000 614.980 1.120 ;
  LAYER metal3 ;
  RECT 613.860 0.000 614.980 1.120 ;
  LAYER metal2 ;
  RECT 613.860 0.000 614.980 1.120 ;
  LAYER metal1 ;
  RECT 613.860 0.000 614.980 1.120 ;
 END
END DI37
PIN DO36
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 608.900 0.000 610.020 1.120 ;
  LAYER metal3 ;
  RECT 608.900 0.000 610.020 1.120 ;
  LAYER metal2 ;
  RECT 608.900 0.000 610.020 1.120 ;
  LAYER metal1 ;
  RECT 608.900 0.000 610.020 1.120 ;
 END
END DO36
PIN DI36
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 600.840 0.000 601.960 1.120 ;
  LAYER metal3 ;
  RECT 600.840 0.000 601.960 1.120 ;
  LAYER metal2 ;
  RECT 600.840 0.000 601.960 1.120 ;
  LAYER metal1 ;
  RECT 600.840 0.000 601.960 1.120 ;
 END
END DI36
PIN DO35
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 595.880 0.000 597.000 1.120 ;
  LAYER metal3 ;
  RECT 595.880 0.000 597.000 1.120 ;
  LAYER metal2 ;
  RECT 595.880 0.000 597.000 1.120 ;
  LAYER metal1 ;
  RECT 595.880 0.000 597.000 1.120 ;
 END
END DO35
PIN DI35
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 587.820 0.000 588.940 1.120 ;
  LAYER metal3 ;
  RECT 587.820 0.000 588.940 1.120 ;
  LAYER metal2 ;
  RECT 587.820 0.000 588.940 1.120 ;
  LAYER metal1 ;
  RECT 587.820 0.000 588.940 1.120 ;
 END
END DI35
PIN DO34
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 582.860 0.000 583.980 1.120 ;
  LAYER metal3 ;
  RECT 582.860 0.000 583.980 1.120 ;
  LAYER metal2 ;
  RECT 582.860 0.000 583.980 1.120 ;
  LAYER metal1 ;
  RECT 582.860 0.000 583.980 1.120 ;
 END
END DO34
PIN DI34
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 574.180 0.000 575.300 1.120 ;
  LAYER metal3 ;
  RECT 574.180 0.000 575.300 1.120 ;
  LAYER metal2 ;
  RECT 574.180 0.000 575.300 1.120 ;
  LAYER metal1 ;
  RECT 574.180 0.000 575.300 1.120 ;
 END
END DI34
PIN DO33
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 566.120 0.000 567.240 1.120 ;
  LAYER metal3 ;
  RECT 566.120 0.000 567.240 1.120 ;
  LAYER metal2 ;
  RECT 566.120 0.000 567.240 1.120 ;
  LAYER metal1 ;
  RECT 566.120 0.000 567.240 1.120 ;
 END
END DO33
PIN DI33
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 557.440 0.000 558.560 1.120 ;
  LAYER metal3 ;
  RECT 557.440 0.000 558.560 1.120 ;
  LAYER metal2 ;
  RECT 557.440 0.000 558.560 1.120 ;
  LAYER metal1 ;
  RECT 557.440 0.000 558.560 1.120 ;
 END
END DI33
PIN DO32
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 552.480 0.000 553.600 1.120 ;
  LAYER metal3 ;
  RECT 552.480 0.000 553.600 1.120 ;
  LAYER metal2 ;
  RECT 552.480 0.000 553.600 1.120 ;
  LAYER metal1 ;
  RECT 552.480 0.000 553.600 1.120 ;
 END
END DO32
PIN DI32
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 544.420 0.000 545.540 1.120 ;
  LAYER metal3 ;
  RECT 544.420 0.000 545.540 1.120 ;
  LAYER metal2 ;
  RECT 544.420 0.000 545.540 1.120 ;
  LAYER metal1 ;
  RECT 544.420 0.000 545.540 1.120 ;
 END
END DI32
PIN DO31
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 539.460 0.000 540.580 1.120 ;
  LAYER metal3 ;
  RECT 539.460 0.000 540.580 1.120 ;
  LAYER metal2 ;
  RECT 539.460 0.000 540.580 1.120 ;
  LAYER metal1 ;
  RECT 539.460 0.000 540.580 1.120 ;
 END
END DO31
PIN DI31
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 530.780 0.000 531.900 1.120 ;
  LAYER metal3 ;
  RECT 530.780 0.000 531.900 1.120 ;
  LAYER metal2 ;
  RECT 530.780 0.000 531.900 1.120 ;
  LAYER metal1 ;
  RECT 530.780 0.000 531.900 1.120 ;
 END
END DI31
PIN DO30
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 525.820 0.000 526.940 1.120 ;
  LAYER metal3 ;
  RECT 525.820 0.000 526.940 1.120 ;
  LAYER metal2 ;
  RECT 525.820 0.000 526.940 1.120 ;
  LAYER metal1 ;
  RECT 525.820 0.000 526.940 1.120 ;
 END
END DO30
PIN DI30
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 517.760 0.000 518.880 1.120 ;
  LAYER metal3 ;
  RECT 517.760 0.000 518.880 1.120 ;
  LAYER metal2 ;
  RECT 517.760 0.000 518.880 1.120 ;
  LAYER metal1 ;
  RECT 517.760 0.000 518.880 1.120 ;
 END
END DI30
PIN DO29
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 509.700 0.000 510.820 1.120 ;
  LAYER metal3 ;
  RECT 509.700 0.000 510.820 1.120 ;
  LAYER metal2 ;
  RECT 509.700 0.000 510.820 1.120 ;
  LAYER metal1 ;
  RECT 509.700 0.000 510.820 1.120 ;
 END
END DO29
PIN DI29
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 501.020 0.000 502.140 1.120 ;
  LAYER metal3 ;
  RECT 501.020 0.000 502.140 1.120 ;
  LAYER metal2 ;
  RECT 501.020 0.000 502.140 1.120 ;
  LAYER metal1 ;
  RECT 501.020 0.000 502.140 1.120 ;
 END
END DI29
PIN DO28
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 496.060 0.000 497.180 1.120 ;
  LAYER metal3 ;
  RECT 496.060 0.000 497.180 1.120 ;
  LAYER metal2 ;
  RECT 496.060 0.000 497.180 1.120 ;
  LAYER metal1 ;
  RECT 496.060 0.000 497.180 1.120 ;
 END
END DO28
PIN DI28
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 488.000 0.000 489.120 1.120 ;
  LAYER metal3 ;
  RECT 488.000 0.000 489.120 1.120 ;
  LAYER metal2 ;
  RECT 488.000 0.000 489.120 1.120 ;
  LAYER metal1 ;
  RECT 488.000 0.000 489.120 1.120 ;
 END
END DI28
PIN DO27
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 483.040 0.000 484.160 1.120 ;
  LAYER metal3 ;
  RECT 483.040 0.000 484.160 1.120 ;
  LAYER metal2 ;
  RECT 483.040 0.000 484.160 1.120 ;
  LAYER metal1 ;
  RECT 483.040 0.000 484.160 1.120 ;
 END
END DO27
PIN DI27
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 474.360 0.000 475.480 1.120 ;
  LAYER metal3 ;
  RECT 474.360 0.000 475.480 1.120 ;
  LAYER metal2 ;
  RECT 474.360 0.000 475.480 1.120 ;
  LAYER metal1 ;
  RECT 474.360 0.000 475.480 1.120 ;
 END
END DI27
PIN DO26
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 469.400 0.000 470.520 1.120 ;
  LAYER metal3 ;
  RECT 469.400 0.000 470.520 1.120 ;
  LAYER metal2 ;
  RECT 469.400 0.000 470.520 1.120 ;
  LAYER metal1 ;
  RECT 469.400 0.000 470.520 1.120 ;
 END
END DO26
PIN DI26
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 461.340 0.000 462.460 1.120 ;
  LAYER metal3 ;
  RECT 461.340 0.000 462.460 1.120 ;
  LAYER metal2 ;
  RECT 461.340 0.000 462.460 1.120 ;
  LAYER metal1 ;
  RECT 461.340 0.000 462.460 1.120 ;
 END
END DI26
PIN DO25
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 452.660 0.000 453.780 1.120 ;
  LAYER metal3 ;
  RECT 452.660 0.000 453.780 1.120 ;
  LAYER metal2 ;
  RECT 452.660 0.000 453.780 1.120 ;
  LAYER metal1 ;
  RECT 452.660 0.000 453.780 1.120 ;
 END
END DO25
PIN DI25
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 444.600 0.000 445.720 1.120 ;
  LAYER metal3 ;
  RECT 444.600 0.000 445.720 1.120 ;
  LAYER metal2 ;
  RECT 444.600 0.000 445.720 1.120 ;
  LAYER metal1 ;
  RECT 444.600 0.000 445.720 1.120 ;
 END
END DI25
PIN DO24
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 439.640 0.000 440.760 1.120 ;
  LAYER metal3 ;
  RECT 439.640 0.000 440.760 1.120 ;
  LAYER metal2 ;
  RECT 439.640 0.000 440.760 1.120 ;
  LAYER metal1 ;
  RECT 439.640 0.000 440.760 1.120 ;
 END
END DO24
PIN DI24
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 430.960 0.000 432.080 1.120 ;
  LAYER metal3 ;
  RECT 430.960 0.000 432.080 1.120 ;
  LAYER metal2 ;
  RECT 430.960 0.000 432.080 1.120 ;
  LAYER metal1 ;
  RECT 430.960 0.000 432.080 1.120 ;
 END
END DI24
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 425.380 0.000 426.500 1.120 ;
  LAYER metal3 ;
  RECT 425.380 0.000 426.500 1.120 ;
  LAYER metal2 ;
  RECT 425.380 0.000 426.500 1.120 ;
  LAYER metal1 ;
  RECT 425.380 0.000 426.500 1.120 ;
 END
END A1
PIN WEB
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 423.520 0.000 424.640 1.120 ;
  LAYER metal3 ;
  RECT 423.520 0.000 424.640 1.120 ;
  LAYER metal2 ;
  RECT 423.520 0.000 424.640 1.120 ;
  LAYER metal1 ;
  RECT 423.520 0.000 424.640 1.120 ;
 END
END WEB
PIN OE
  DIRECTION INPUT ;
  CAPACITANCE 0.033 ;
 PORT
  LAYER metal4 ;
  RECT 419.180 0.000 420.300 1.120 ;
  LAYER metal3 ;
  RECT 419.180 0.000 420.300 1.120 ;
  LAYER metal2 ;
  RECT 419.180 0.000 420.300 1.120 ;
  LAYER metal1 ;
  RECT 419.180 0.000 420.300 1.120 ;
 END
END OE
PIN CS
  DIRECTION INPUT ;
  CAPACITANCE 0.123 ;
 PORT
  LAYER metal4 ;
  RECT 417.320 0.000 418.440 1.120 ;
  LAYER metal3 ;
  RECT 417.320 0.000 418.440 1.120 ;
  LAYER metal2 ;
  RECT 417.320 0.000 418.440 1.120 ;
  LAYER metal1 ;
  RECT 417.320 0.000 418.440 1.120 ;
 END
END CS
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 395.620 0.000 396.740 1.120 ;
  LAYER metal3 ;
  RECT 395.620 0.000 396.740 1.120 ;
  LAYER metal2 ;
  RECT 395.620 0.000 396.740 1.120 ;
  LAYER metal1 ;
  RECT 395.620 0.000 396.740 1.120 ;
 END
END A2
PIN CK
  DIRECTION INPUT ;
  CAPACITANCE 0.063 ;
 PORT
  LAYER metal4 ;
  RECT 392.520 0.000 393.640 1.120 ;
  LAYER metal3 ;
  RECT 392.520 0.000 393.640 1.120 ;
  LAYER metal2 ;
  RECT 392.520 0.000 393.640 1.120 ;
  LAYER metal1 ;
  RECT 392.520 0.000 393.640 1.120 ;
 END
END CK
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 390.040 0.000 391.160 1.120 ;
  LAYER metal3 ;
  RECT 390.040 0.000 391.160 1.120 ;
  LAYER metal2 ;
  RECT 390.040 0.000 391.160 1.120 ;
  LAYER metal1 ;
  RECT 390.040 0.000 391.160 1.120 ;
 END
END A0
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 385.700 0.000 386.820 1.120 ;
  LAYER metal3 ;
  RECT 385.700 0.000 386.820 1.120 ;
  LAYER metal2 ;
  RECT 385.700 0.000 386.820 1.120 ;
  LAYER metal1 ;
  RECT 385.700 0.000 386.820 1.120 ;
 END
END A3
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 378.260 0.000 379.380 1.120 ;
  LAYER metal3 ;
  RECT 378.260 0.000 379.380 1.120 ;
  LAYER metal2 ;
  RECT 378.260 0.000 379.380 1.120 ;
  LAYER metal1 ;
  RECT 378.260 0.000 379.380 1.120 ;
 END
END A4
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 375.160 0.000 376.280 1.120 ;
  LAYER metal3 ;
  RECT 375.160 0.000 376.280 1.120 ;
  LAYER metal2 ;
  RECT 375.160 0.000 376.280 1.120 ;
  LAYER metal1 ;
  RECT 375.160 0.000 376.280 1.120 ;
 END
END A5
PIN A6
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 367.720 0.000 368.840 1.120 ;
  LAYER metal3 ;
  RECT 367.720 0.000 368.840 1.120 ;
  LAYER metal2 ;
  RECT 367.720 0.000 368.840 1.120 ;
  LAYER metal1 ;
  RECT 367.720 0.000 368.840 1.120 ;
 END
END A6
PIN A7
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 364.620 0.000 365.740 1.120 ;
  LAYER metal3 ;
  RECT 364.620 0.000 365.740 1.120 ;
  LAYER metal2 ;
  RECT 364.620 0.000 365.740 1.120 ;
  LAYER metal1 ;
  RECT 364.620 0.000 365.740 1.120 ;
 END
END A7
PIN A8
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 357.180 0.000 358.300 1.120 ;
  LAYER metal3 ;
  RECT 357.180 0.000 358.300 1.120 ;
  LAYER metal2 ;
  RECT 357.180 0.000 358.300 1.120 ;
  LAYER metal1 ;
  RECT 357.180 0.000 358.300 1.120 ;
 END
END A8
PIN DO23
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 346.020 0.000 347.140 1.120 ;
  LAYER metal3 ;
  RECT 346.020 0.000 347.140 1.120 ;
  LAYER metal2 ;
  RECT 346.020 0.000 347.140 1.120 ;
  LAYER metal1 ;
  RECT 346.020 0.000 347.140 1.120 ;
 END
END DO23
PIN DI23
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 337.340 0.000 338.460 1.120 ;
  LAYER metal3 ;
  RECT 337.340 0.000 338.460 1.120 ;
  LAYER metal2 ;
  RECT 337.340 0.000 338.460 1.120 ;
  LAYER metal1 ;
  RECT 337.340 0.000 338.460 1.120 ;
 END
END DI23
PIN DO22
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 332.380 0.000 333.500 1.120 ;
  LAYER metal3 ;
  RECT 332.380 0.000 333.500 1.120 ;
  LAYER metal2 ;
  RECT 332.380 0.000 333.500 1.120 ;
  LAYER metal1 ;
  RECT 332.380 0.000 333.500 1.120 ;
 END
END DO22
PIN DI22
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 324.320 0.000 325.440 1.120 ;
  LAYER metal3 ;
  RECT 324.320 0.000 325.440 1.120 ;
  LAYER metal2 ;
  RECT 324.320 0.000 325.440 1.120 ;
  LAYER metal1 ;
  RECT 324.320 0.000 325.440 1.120 ;
 END
END DI22
PIN DO21
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 316.260 0.000 317.380 1.120 ;
  LAYER metal3 ;
  RECT 316.260 0.000 317.380 1.120 ;
  LAYER metal2 ;
  RECT 316.260 0.000 317.380 1.120 ;
  LAYER metal1 ;
  RECT 316.260 0.000 317.380 1.120 ;
 END
END DO21
PIN DI21
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 307.580 0.000 308.700 1.120 ;
  LAYER metal3 ;
  RECT 307.580 0.000 308.700 1.120 ;
  LAYER metal2 ;
  RECT 307.580 0.000 308.700 1.120 ;
  LAYER metal1 ;
  RECT 307.580 0.000 308.700 1.120 ;
 END
END DI21
PIN DO20
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 302.620 0.000 303.740 1.120 ;
  LAYER metal3 ;
  RECT 302.620 0.000 303.740 1.120 ;
  LAYER metal2 ;
  RECT 302.620 0.000 303.740 1.120 ;
  LAYER metal1 ;
  RECT 302.620 0.000 303.740 1.120 ;
 END
END DO20
PIN DI20
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 294.560 0.000 295.680 1.120 ;
  LAYER metal3 ;
  RECT 294.560 0.000 295.680 1.120 ;
  LAYER metal2 ;
  RECT 294.560 0.000 295.680 1.120 ;
  LAYER metal1 ;
  RECT 294.560 0.000 295.680 1.120 ;
 END
END DI20
PIN DO19
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 289.600 0.000 290.720 1.120 ;
  LAYER metal3 ;
  RECT 289.600 0.000 290.720 1.120 ;
  LAYER metal2 ;
  RECT 289.600 0.000 290.720 1.120 ;
  LAYER metal1 ;
  RECT 289.600 0.000 290.720 1.120 ;
 END
END DO19
PIN DI19
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 280.920 0.000 282.040 1.120 ;
  LAYER metal3 ;
  RECT 280.920 0.000 282.040 1.120 ;
  LAYER metal2 ;
  RECT 280.920 0.000 282.040 1.120 ;
  LAYER metal1 ;
  RECT 280.920 0.000 282.040 1.120 ;
 END
END DI19
PIN DO18
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 275.960 0.000 277.080 1.120 ;
  LAYER metal3 ;
  RECT 275.960 0.000 277.080 1.120 ;
  LAYER metal2 ;
  RECT 275.960 0.000 277.080 1.120 ;
  LAYER metal1 ;
  RECT 275.960 0.000 277.080 1.120 ;
 END
END DO18
PIN DI18
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal3 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal2 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal1 ;
  RECT 267.900 0.000 269.020 1.120 ;
 END
END DI18
PIN DO17
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER metal3 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER metal2 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER metal1 ;
  RECT 259.220 0.000 260.340 1.120 ;
 END
END DO17
PIN DI17
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER metal3 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER metal2 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER metal1 ;
  RECT 251.160 0.000 252.280 1.120 ;
 END
END DI17
PIN DO16
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER metal3 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER metal2 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER metal1 ;
  RECT 246.200 0.000 247.320 1.120 ;
 END
END DO16
PIN DI16
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER metal3 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER metal2 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER metal1 ;
  RECT 237.520 0.000 238.640 1.120 ;
 END
END DI16
PIN DO15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER metal3 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER metal2 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER metal1 ;
  RECT 233.180 0.000 234.300 1.120 ;
 END
END DO15
PIN DI15
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER metal3 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER metal2 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER metal1 ;
  RECT 224.500 0.000 225.620 1.120 ;
 END
END DI15
PIN DO14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER metal3 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER metal2 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER metal1 ;
  RECT 219.540 0.000 220.660 1.120 ;
 END
END DO14
PIN DI14
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER metal3 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER metal2 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER metal1 ;
  RECT 211.480 0.000 212.600 1.120 ;
 END
END DI14
PIN DO13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER metal3 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER metal2 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER metal1 ;
  RECT 202.800 0.000 203.920 1.120 ;
 END
END DO13
PIN DI13
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER metal3 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER metal2 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER metal1 ;
  RECT 194.740 0.000 195.860 1.120 ;
 END
END DI13
PIN DO12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER metal3 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER metal2 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER metal1 ;
  RECT 189.780 0.000 190.900 1.120 ;
 END
END DO12
PIN DI12
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER metal3 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER metal2 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER metal1 ;
  RECT 181.100 0.000 182.220 1.120 ;
 END
END DI12
PIN DO11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER metal3 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER metal2 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER metal1 ;
  RECT 176.140 0.000 177.260 1.120 ;
 END
END DO11
PIN DI11
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER metal3 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER metal2 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER metal1 ;
  RECT 168.080 0.000 169.200 1.120 ;
 END
END DI11
PIN DO10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER metal3 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER metal2 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER metal1 ;
  RECT 163.120 0.000 164.240 1.120 ;
 END
END DO10
PIN DI10
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER metal3 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER metal2 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER metal1 ;
  RECT 154.440 0.000 155.560 1.120 ;
 END
END DI10
PIN DO9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER metal3 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER metal2 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER metal1 ;
  RECT 146.380 0.000 147.500 1.120 ;
 END
END DO9
PIN DI9
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER metal3 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER metal2 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER metal1 ;
  RECT 137.700 0.000 138.820 1.120 ;
 END
END DI9
PIN DO8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER metal3 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER metal2 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER metal1 ;
  RECT 133.360 0.000 134.480 1.120 ;
 END
END DO8
PIN DI8
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER metal3 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER metal2 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER metal1 ;
  RECT 124.680 0.000 125.800 1.120 ;
 END
END DI8
PIN DO7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER metal3 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER metal2 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER metal1 ;
  RECT 119.720 0.000 120.840 1.120 ;
 END
END DO7
PIN DI7
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER metal3 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER metal2 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER metal1 ;
  RECT 111.660 0.000 112.780 1.120 ;
 END
END DI7
PIN DO6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal3 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal2 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal1 ;
  RECT 106.700 0.000 107.820 1.120 ;
 END
END DO6
PIN DI6
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER metal3 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER metal2 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER metal1 ;
  RECT 98.020 0.000 99.140 1.120 ;
 END
END DI6
PIN DO5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER metal3 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER metal2 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER metal1 ;
  RECT 89.960 0.000 91.080 1.120 ;
 END
END DO5
PIN DI5
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER metal3 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER metal2 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER metal1 ;
  RECT 81.280 0.000 82.400 1.120 ;
 END
END DI5
PIN DO4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER metal3 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER metal2 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER metal1 ;
  RECT 76.320 0.000 77.440 1.120 ;
 END
END DO4
PIN DI4
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER metal3 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER metal2 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER metal1 ;
  RECT 68.260 0.000 69.380 1.120 ;
 END
END DI4
PIN DO3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER metal3 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER metal2 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER metal1 ;
  RECT 63.300 0.000 64.420 1.120 ;
 END
END DO3
PIN DI3
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER metal3 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER metal2 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER metal1 ;
  RECT 54.620 0.000 55.740 1.120 ;
 END
END DI3
PIN DO2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER metal3 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER metal2 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER metal1 ;
  RECT 50.280 0.000 51.400 1.120 ;
 END
END DO2
PIN DI2
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER metal3 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER metal2 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER metal1 ;
  RECT 41.600 0.000 42.720 1.120 ;
 END
END DI2
PIN DO1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal3 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal2 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal1 ;
  RECT 33.540 0.000 34.660 1.120 ;
 END
END DO1
PIN DI1
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal3 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal2 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal1 ;
  RECT 24.860 0.000 25.980 1.120 ;
 END
END DI1
PIN DO0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal3 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal2 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal1 ;
  RECT 19.900 0.000 21.020 1.120 ;
 END
END DO0
PIN DI0
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal3 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal2 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal1 ;
  RECT 11.840 0.000 12.960 1.120 ;
 END
END DI0
OBS
  LAYER metal1 SPACING 0.280 ;
  RECT 0.000 0.140 778.720 225.680 ;
  LAYER metal2 SPACING 0.320 ;
  RECT 0.000 0.140 778.720 225.680 ;
  LAYER metal3 SPACING 0.320 ;
  RECT 0.000 0.140 778.720 225.680 ;
  LAYER metal4 SPACING 0.600 ;
  RECT 0.000 0.140 778.720 225.680 ;
  LAYER via ;
  RECT 0.000 0.140 778.720 225.680 ;
  LAYER via2 ;
  RECT 0.000 0.140 778.720 225.680 ;
  LAYER via3 ;
  RECT 0.000 0.140 778.720 225.680 ;
END
END SUMA180_288X48X1BM1
END LIBRARY



